module get_tse_data 
   (
		output 		[7:0] gmac_tx_data_1_out,
		output 		gmac_tx_dvld_1_out,
		output 		gmac_tx_ack_1_out,
		  
		input 		[7:0] gmac_rx_data_1_in,
		input 		gmac_rx_dvld_1_in,
		input 		gmac_rx_frame_error_1_in, 

      // core clock
      input        core_clk_int,

      // misc
      input        reset    

   );
	
	
	
	
	
	endmodule