//
//	8192 bytes, 32bit interface

`timescale 1ns/1ps


module bb_ram(clk, addr, data_in, data_out, we, en, reset);
input clk;
input [12:2] addr;
input [31:0] data_in;
output [31:0] data_out;
input [3:0] we;
input en;
input reset;

wire [3:0] dip;

RAMB16_S9 ram0(

        .DO     (data_out[7:0]),
	.DOP    (),
	.ADDR   (addr[12:2]),
	.CLK    (clk),
	.DI     (data_in[7:0]),
	.DIP    (dip[0]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[0])

);

defparam ram0.INIT_00 = 256'h0505050505050505050505040303030303030303020202020202020201010101;
defparam ram0.INIT_01 = 256'h0505050505050505050505050505050505050505050505050505050505050505;
defparam ram0.INIT_02 = 256'h0707070707070707070707070706060605050505050505050505050505050505;
defparam ram0.INIT_03 = 256'h0909090909080807070707070707070707070707070707070707070707070707;
defparam ram0.INIT_04 = 256'h0D0D0D0C0C0C0C0C0C0C0C0C0C0C0B0B0A0A0A0A0A0A0A0A0A0A0A0A0A0A0A09;
defparam ram0.INIT_05 = 256'h00000000101010101010100F0F0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0D0D;
defparam ram0.INIT_06 = 256'h0000000000000000000000000000;
defparam ram0.INIT_07 = 256'h0000000000000000000000000000;
defparam ram0.INIT_08 = 256'h0000000000000000000000000000;
defparam ram0.INIT_09 = 256'h0000000000000000000000000000;
defparam ram0.INIT_0A = 256'h0000000000000000000000000000;
defparam ram0.INIT_0B = 256'h0000000000000000000000000000;
defparam ram0.INIT_0C = 256'h0000000000000000000000000000;
defparam ram0.INIT_0D = 256'h0000000000000000000000000000;
defparam ram0.INIT_0E = 256'h0000000000000000000000000000;
defparam ram0.INIT_0F = 256'h0000000000000000000000000000;
defparam ram0.INIT_10 = 256'h0000000000000000000000000000;
defparam ram0.INIT_11 = 256'h0000000000000000000000000000;
defparam ram0.INIT_12 = 256'h0000000000000000000000000000;
defparam ram0.INIT_13 = 256'h0000000000000000000000000000;
defparam ram0.INIT_14 = 256'h0000000000000000000000000000;
defparam ram0.INIT_15 = 256'h0000000000000000000000000000;
defparam ram0.INIT_16 = 256'h0000000000000000000000000000;
defparam ram0.INIT_17 = 256'h0000000000000000000000000000;
defparam ram0.INIT_18 = 256'h0000000000000000000000000000;
defparam ram0.INIT_19 = 256'h0000000000000000000000000000;
defparam ram0.INIT_1A = 256'h0000000000000000000000000000;
defparam ram0.INIT_1B = 256'h0000000000000000000000000000;
defparam ram0.INIT_1C = 256'h0000000000000000000000000000;
defparam ram0.INIT_1D = 256'h0000000000000000000000000000;
defparam ram0.INIT_1E = 256'h0000000000000000000000000000;
defparam ram0.INIT_1F = 256'h0000000000000000000000000000;
defparam ram0.INIT_20 = 256'h0000000000000000000000000000;
defparam ram0.INIT_21 = 256'h0000000000000000000000000000;
defparam ram0.INIT_22 = 256'h0000000000000000000000000000;
defparam ram0.INIT_23 = 256'h0000000000000000000000000000;
defparam ram0.INIT_24 = 256'h0000000000000000000000000000;
defparam ram0.INIT_25 = 256'h0000000000000000000000000000;
defparam ram0.INIT_26 = 256'h0000000000000000000000000000;
defparam ram0.INIT_27 = 256'h0000000000000000000000000000;
defparam ram0.INIT_28 = 256'h0000000000000000000000000000;
defparam ram0.INIT_29 = 256'h0000000000000000000000000000;
defparam ram0.INIT_2A = 256'h0000000000000000000000000000;
defparam ram0.INIT_2B = 256'h0000000000000000000000000000;
defparam ram0.INIT_2C = 256'h0000000000000000000000000000;
defparam ram0.INIT_2D = 256'h0000000000000000000000000000;
defparam ram0.INIT_2E = 256'h0000000000000000000000000000;
defparam ram0.INIT_2F = 256'h0000000000000000000000000000;
defparam ram0.INIT_30 = 256'h0000000000000000000000000000;
defparam ram0.INIT_31 = 256'h0000000000000000000000000000;
defparam ram0.INIT_32 = 256'h0000000000000000000000000000;
defparam ram0.INIT_33 = 256'h0000000000000000000000000000;
defparam ram0.INIT_34 = 256'h0000000000000000000000000000;
defparam ram0.INIT_35 = 256'h0000000000000000000000000000;
defparam ram0.INIT_36 = 256'h0000000000000000000000000000;
defparam ram0.INIT_37 = 256'h0000000000000000000000000000;
defparam ram0.INIT_38 = 256'h0000000000000000000000000000;
defparam ram0.INIT_39 = 256'h0000000000000000000000000000;
defparam ram0.INIT_3A = 256'h0000000000000000000000000000;
defparam ram0.INIT_3B = 256'h0000000000000000000000000000;
defparam ram0.INIT_3C = 256'h0000000000000000000000000000;
defparam ram0.INIT_3D = 256'h0000000000000000000000000000;
defparam ram0.INIT_3E = 256'h0000000000000000000000000000;
defparam ram0.INIT_3F = 256'h0000000000000000000000000000;


RAMB16_S9 ram1(

        .DO     (data_out[15:8]),
	.DOP    (),
	.ADDR   (addr[12:2]),
	.CLK    (clk),
	.DI     (data_in[15:8]),
	.DIP    (dip[1]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[1])

);

defparam ram1.INIT_00 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_01 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_02 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_03 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_04 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_05 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_06 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_07 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_08 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_09 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0A = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0B = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0C = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0D = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0E = 256'h00000000000000000000000000000000;
defparam ram1.INIT_0F = 256'h00000000000000000000000000000000;
defparam ram1.INIT_10 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_11 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_12 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_13 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_14 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_15 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_16 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_17 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_18 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_19 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1A = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1B = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1C = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1D = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1E = 256'h00000000000000000000000000000000;
defparam ram1.INIT_1F = 256'h00000000000000000000000000000000;
defparam ram1.INIT_20 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_21 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_22 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_23 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_24 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_25 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_26 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_27 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_28 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_29 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2A = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2B = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2C = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2D = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2E = 256'h00000000000000000000000000000000;
defparam ram1.INIT_2F = 256'h00000000000000000000000000000000;
defparam ram1.INIT_30 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_31 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_32 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_33 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_34 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_35 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_36 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_37 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_38 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_39 = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3A = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3B = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3C = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3D = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3E = 256'h00000000000000000000000000000000;
defparam ram1.INIT_3F = 256'h00000000000000000000000000000000;


RAMB16_S9 ram2(

        .DO     (data_out[23:16]),
	.DOP    (),
	.ADDR   (addr[12:2]),
	.CLK    (clk),
	.DI     (data_in[23:16]),
	.DIP    (dip[2]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[2])

);
defparam ram2.INIT_00 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_01 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_02 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_03 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_04 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_05 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_06 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_07 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_08 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_09 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0A = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0B = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0C = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0D = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0E = 256'h00000000000000000000000000000000;
defparam ram2.INIT_0F = 256'h00000000000000000000000000000000;
defparam ram2.INIT_10 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_11 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_12 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_13 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_14 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_15 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_16 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_17 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_18 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_19 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1A = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1B = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1C = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1D = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1E = 256'h00000000000000000000000000000000;
defparam ram2.INIT_1F = 256'h00000000000000000000000000000000;
defparam ram2.INIT_20 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_21 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_22 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_23 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_24 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_25 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_26 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_27 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_28 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_29 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2A = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2B = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2C = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2D = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2E = 256'h00000000000000000000000000000000;
defparam ram2.INIT_2F = 256'h00000000000000000000000000000000;
defparam ram2.INIT_30 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_31 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_32 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_33 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_34 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_35 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_36 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_37 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_38 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_39 = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3A = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3B = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3C = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3D = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3E = 256'h00000000000000000000000000000000;
defparam ram2.INIT_3F = 256'h00000000000000000000000000000000;



RAMB16_S9 ram3(

        .DO     (data_out[31:24]),
	.DOP    (),
	.ADDR   (addr[12:2]),
	.CLK    (clk),
	.DI     (data_in[31:24]),
	.DIP    (dip[3]),
	.EN     (en),
	.SSR    (reset),
	.WE     (we[3])

);

defparam ram3.INIT_00 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_01 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_02 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_03 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_04 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_05 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_06 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_07 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_08 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_09 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0A = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0B = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0C = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0D = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0E = 256'h00000000000000000000000000000000;
defparam ram3.INIT_0F = 256'h00000000000000000000000000000000;
defparam ram3.INIT_10 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_11 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_12 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_13 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_14 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_15 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_16 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_17 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_18 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_19 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1A = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1B = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1C = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1D = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1E = 256'h00000000000000000000000000000000;
defparam ram3.INIT_1F = 256'h00000000000000000000000000000000;
defparam ram3.INIT_20 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_21 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_22 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_23 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_24 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_25 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_26 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_27 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_28 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_29 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2A = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2B = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2C = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2D = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2E = 256'h00000000000000000000000000000000;
defparam ram3.INIT_2F = 256'h00000000000000000000000000000000;
defparam ram3.INIT_30 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_31 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_32 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_33 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_34 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_35 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_36 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_37 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_38 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_39 = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3A = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3B = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3C = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3D = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3E = 256'h00000000000000000000000000000000;
defparam ram3.INIT_3F = 256'h00000000000000000000000000000000;

endmodule
