library verilog;
use verilog.vl_types.all;
entity flow_classification is
    generic(
        PRO_IDLE        : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        PRO_FIND1       : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        PRO_FIND2       : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        PRO_FIND3       : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        PRO_FIND4       : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        FC_IDLE         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        FC_LOOKUP_ROUTE : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        FC_REQ          : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        FC_ACK          : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        FC_TX           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        FC_CANCEL_REQ   : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        FC_WAIT_ACK     : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1)
    );
    port(
        out_data0       : out    vl_logic_vector(63 downto 0);
        out_pkt_route0  : out    vl_logic_vector(23 downto 0);
        out_wr0         : out    vl_logic;
        out_req0        : out    vl_logic;
        out_ack0        : in     vl_logic;
        out_bypass0     : out    vl_logic;
        out_protocol0   : out    vl_logic;
        out_data1       : out    vl_logic_vector(63 downto 0);
        out_pkt_route1  : out    vl_logic_vector(23 downto 0);
        out_wr1         : out    vl_logic;
        out_req1        : out    vl_logic;
        out_ack1        : in     vl_logic;
        out_bypass1     : out    vl_logic;
        out_protocol1   : out    vl_logic;
        out_data2       : out    vl_logic_vector(63 downto 0);
        out_pkt_route2  : out    vl_logic_vector(23 downto 0);
        out_wr2         : out    vl_logic;
        out_req2        : out    vl_logic;
        out_ack2        : in     vl_logic;
        out_bypass2     : out    vl_logic;
        out_protocol2   : out    vl_logic;
        out_data3       : out    vl_logic_vector(63 downto 0);
        out_pkt_route3  : out    vl_logic_vector(23 downto 0);
        out_wr3         : out    vl_logic;
        out_req3        : out    vl_logic;
        out_ack3        : in     vl_logic;
        out_bypass3     : out    vl_logic;
        out_protocol3   : out    vl_logic;
        in_data         : in     vl_logic_vector(63 downto 0);
        in_ctrl         : in     vl_logic_vector(7 downto 0);
        in_wr           : in     vl_logic;
        in_rdy          : out    vl_logic;
        reg_req_in      : in     vl_logic;
        reg_ack_in      : in     vl_logic;
        reg_rd_wr_L_in  : in     vl_logic;
        reg_addr_in     : in     vl_logic_vector(22 downto 0);
        reg_data_in     : in     vl_logic_vector(31 downto 0);
        reg_src_in      : in     vl_logic_vector(1 downto 0);
        reg_req_out     : out    vl_logic;
        reg_ack_out     : out    vl_logic;
        reg_rd_wr_L_out : out    vl_logic;
        reg_addr_out    : out    vl_logic_vector(22 downto 0);
        reg_data_out    : out    vl_logic_vector(31 downto 0);
        reg_src_out     : out    vl_logic_vector(1 downto 0);
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        protocol_signal : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of PRO_IDLE : constant is 1;
    attribute mti_svvh_generic_type of PRO_FIND1 : constant is 1;
    attribute mti_svvh_generic_type of PRO_FIND2 : constant is 1;
    attribute mti_svvh_generic_type of PRO_FIND3 : constant is 1;
    attribute mti_svvh_generic_type of PRO_FIND4 : constant is 1;
    attribute mti_svvh_generic_type of FC_IDLE : constant is 1;
    attribute mti_svvh_generic_type of FC_LOOKUP_ROUTE : constant is 1;
    attribute mti_svvh_generic_type of FC_REQ : constant is 1;
    attribute mti_svvh_generic_type of FC_ACK : constant is 1;
    attribute mti_svvh_generic_type of FC_TX : constant is 1;
    attribute mti_svvh_generic_type of FC_CANCEL_REQ : constant is 1;
    attribute mti_svvh_generic_type of FC_WAIT_ACK : constant is 1;
end flow_classification;
