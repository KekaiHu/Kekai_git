library verilog;
use verilog.vl_types.all;
entity unused_reg is
    generic(
        REG_ADDR_WIDTH  : integer := 5
    );
    port(
        reg_req         : in     vl_logic;
        reg_ack         : out    vl_logic;
        reg_rd_wr_L     : in     vl_logic;
        reg_addr        : in     vl_logic_vector;
        reg_rd_data     : out    vl_logic_vector(31 downto 0);
        reg_wr_data     : in     vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of REG_ADDR_WIDTH : constant is 1;
end unused_reg;
