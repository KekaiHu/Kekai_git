library verilog;
use verilog.vl_types.all;
entity fallthrough_small_fifo_tester is
end fallthrough_small_fifo_tester;
