library verilog;
use verilog.vl_types.all;
entity ppu is
    generic(
        SP_IDLE         : vl_logic := Hi0;
        SP_PROC         : vl_logic := Hi1
    );
    port(
        clk             : in     vl_logic;
        core_sp_clk     : in     vl_logic;
        reset           : in     vl_logic;
        TRIG_IS         : out    vl_logic_vector(239 downto 0);
        TRIG_OS         : out    vl_logic_vector(239 downto 0);
        in_data0        : in     vl_logic_vector(63 downto 0);
        in_pkt_route0   : in     vl_logic_vector(23 downto 0);
        in_wr0          : in     vl_logic;
        in_req0         : in     vl_logic;
        in_ack0         : out    vl_logic;
        in_bypass0      : in     vl_logic;
        in_data1        : in     vl_logic_vector(63 downto 0);
        in_pkt_route1   : in     vl_logic_vector(23 downto 0);
        in_wr1          : in     vl_logic;
        in_req1         : in     vl_logic;
        in_ack1         : out    vl_logic;
        in_bypass1      : in     vl_logic;
        in_protocol1    : in     vl_logic;
        in_data2        : in     vl_logic_vector(63 downto 0);
        in_pkt_route2   : in     vl_logic_vector(23 downto 0);
        in_wr2          : in     vl_logic;
        in_req2         : in     vl_logic;
        in_ack2         : out    vl_logic;
        in_bypass2      : in     vl_logic;
        in_data3        : in     vl_logic_vector(63 downto 0);
        in_pkt_route3   : in     vl_logic_vector(23 downto 0);
        in_wr3          : in     vl_logic;
        in_req3         : in     vl_logic;
        in_ack3         : out    vl_logic;
        in_bypass3      : in     vl_logic;
        out_data0       : out    vl_logic_vector(63 downto 0);
        out_pkt_route0  : out    vl_logic_vector(23 downto 0);
        out_wr0         : out    vl_logic;
        out_req0        : out    vl_logic;
        out_ack0        : in     vl_logic;
        out_bop0        : out    vl_logic;
        out_eop0        : out    vl_logic;
        out_rdy0        : in     vl_logic;
        out_bypass0     : out    vl_logic;
        out_data1       : out    vl_logic_vector(63 downto 0);
        out_pkt_route1  : out    vl_logic_vector(23 downto 0);
        out_wr1         : out    vl_logic;
        out_req1        : out    vl_logic;
        out_ack1        : in     vl_logic;
        out_bop1        : out    vl_logic;
        out_eop1        : out    vl_logic;
        out_rdy1        : in     vl_logic;
        out_bypass1     : out    vl_logic;
        out_data2       : out    vl_logic_vector(63 downto 0);
        out_pkt_route2  : out    vl_logic_vector(23 downto 0);
        out_wr2         : out    vl_logic;
        out_req2        : out    vl_logic;
        out_ack2        : in     vl_logic;
        out_bop2        : out    vl_logic;
        out_eop2        : out    vl_logic;
        out_rdy2        : in     vl_logic;
        out_bypass2     : out    vl_logic;
        out_data3       : out    vl_logic_vector(63 downto 0);
        out_pkt_route3  : out    vl_logic_vector(23 downto 0);
        out_wr3         : out    vl_logic;
        out_req3        : out    vl_logic;
        out_ack3        : in     vl_logic;
        out_bop3        : out    vl_logic;
        out_eop3        : out    vl_logic;
        out_rdy3        : in     vl_logic;
        out_bypass3     : out    vl_logic;
        cam_we          : in     vl_logic;
        cam_wr_addr     : in     vl_logic_vector(3 downto 0);
        cam_din         : in     vl_logic_vector(31 downto 0);
        cam_wr_ack      : out    vl_logic;
        out_four_bit_hash: out    vl_logic_vector(3 downto 0);
        out_new_inst_signal: out    vl_logic;
        in_packet_drop_signal: in     vl_logic;
        out_ack_reset   : in     vl_logic;
        out_processor_reset_seq: out    vl_logic;
        out_sp_pkt_done : out    vl_logic;
        out_sp_interrupt_wire: out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SP_IDLE : constant is 1;
    attribute mti_svvh_generic_type of SP_PROC : constant is 1;
end ppu;
