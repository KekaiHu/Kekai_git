library verilog;
use verilog.vl_types.all;
entity out_switch is
    generic(
        OS_IDLE         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        OS_LOOKUP_BUFF  : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        OS_PORT_REQ     : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        OS_TX           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        OS_CANCEL       : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1)
    );
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        TRIG0           : out    vl_logic_vector(239 downto 0);
        pb_out_data0    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route0: in     vl_logic_vector(23 downto 0);
        pb_out_wr0      : in     vl_logic;
        pb_out_req0     : in     vl_logic;
        pb_out_ack0     : out    vl_logic;
        pb_out_neighbor0: in     vl_logic_vector(1 downto 0);
        pb_out_bop0     : in     vl_logic;
        pb_out_eop0     : in     vl_logic;
        pb_out_rdy0     : out    vl_logic;
        pb_out_bypass0  : in     vl_logic;
        pb_out_data1    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route1: in     vl_logic_vector(23 downto 0);
        pb_out_wr1      : in     vl_logic;
        pb_out_req1     : in     vl_logic;
        pb_out_ack1     : out    vl_logic;
        pb_out_neighbor1: in     vl_logic_vector(1 downto 0);
        pb_out_bop1     : in     vl_logic;
        pb_out_eop1     : in     vl_logic;
        pb_out_rdy1     : out    vl_logic;
        pb_out_bypass1  : in     vl_logic;
        pb_out_data2    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route2: in     vl_logic_vector(23 downto 0);
        pb_out_wr2      : in     vl_logic;
        pb_out_req2     : in     vl_logic;
        pb_out_ack2     : out    vl_logic;
        pb_out_neighbor2: in     vl_logic_vector(1 downto 0);
        pb_out_bop2     : in     vl_logic;
        pb_out_eop2     : in     vl_logic;
        pb_out_rdy2     : out    vl_logic;
        pb_out_bypass2  : in     vl_logic;
        pb_out_data3    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route3: in     vl_logic_vector(23 downto 0);
        pb_out_wr3      : in     vl_logic;
        pb_out_req3     : in     vl_logic;
        pb_out_ack3     : out    vl_logic;
        pb_out_neighbor3: in     vl_logic_vector(1 downto 0);
        pb_out_bop3     : in     vl_logic;
        pb_out_eop3     : in     vl_logic;
        pb_out_rdy3     : out    vl_logic;
        pb_out_bypass3  : in     vl_logic;
        pb_out_data4    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route4: in     vl_logic_vector(23 downto 0);
        pb_out_wr4      : in     vl_logic;
        pb_out_req4     : in     vl_logic;
        pb_out_ack4     : out    vl_logic;
        pb_out_neighbor4: in     vl_logic_vector(1 downto 0);
        pb_out_bop4     : in     vl_logic;
        pb_out_eop4     : in     vl_logic;
        pb_out_rdy4     : out    vl_logic;
        pb_out_bypass4  : in     vl_logic;
        pb_out_data5    : in     vl_logic_vector(63 downto 0);
        pb_out_pkt_route5: in     vl_logic_vector(23 downto 0);
        pb_out_wr5      : in     vl_logic;
        pb_out_req5     : in     vl_logic;
        pb_out_ack5     : out    vl_logic;
        pb_out_neighbor5: in     vl_logic_vector(1 downto 0);
        pb_out_bop5     : in     vl_logic;
        pb_out_eop5     : in     vl_logic;
        pb_out_rdy5     : out    vl_logic;
        pb_out_bypass5  : in     vl_logic;
        out_data0       : out    vl_logic_vector(63 downto 0);
        out_pkt_route0  : out    vl_logic_vector(23 downto 0);
        out_wr0         : out    vl_logic;
        out_req0        : out    vl_logic;
        out_ack0        : in     vl_logic;
        out_bop0        : out    vl_logic;
        out_eop0        : out    vl_logic;
        out_rdy0        : in     vl_logic;
        out_bypass0     : out    vl_logic;
        out_data1       : out    vl_logic_vector(63 downto 0);
        out_pkt_route1  : out    vl_logic_vector(23 downto 0);
        out_wr1         : out    vl_logic;
        out_req1        : out    vl_logic;
        out_ack1        : in     vl_logic;
        out_bop1        : out    vl_logic;
        out_eop1        : out    vl_logic;
        out_rdy1        : in     vl_logic;
        out_bypass1     : out    vl_logic;
        out_data2       : out    vl_logic_vector(63 downto 0);
        out_pkt_route2  : out    vl_logic_vector(23 downto 0);
        out_wr2         : out    vl_logic;
        out_req2        : out    vl_logic;
        out_ack2        : in     vl_logic;
        out_bop2        : out    vl_logic;
        out_eop2        : out    vl_logic;
        out_rdy2        : in     vl_logic;
        out_bypass2     : out    vl_logic;
        out_data3       : out    vl_logic_vector(63 downto 0);
        out_pkt_route3  : out    vl_logic_vector(23 downto 0);
        out_wr3         : out    vl_logic;
        out_req3        : out    vl_logic;
        out_ack3        : in     vl_logic;
        out_bop3        : out    vl_logic;
        out_eop3        : out    vl_logic;
        out_rdy3        : in     vl_logic;
        out_bypass3     : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of OS_IDLE : constant is 1;
    attribute mti_svvh_generic_type of OS_LOOKUP_BUFF : constant is 1;
    attribute mti_svvh_generic_type of OS_PORT_REQ : constant is 1;
    attribute mti_svvh_generic_type of OS_TX : constant is 1;
    attribute mti_svvh_generic_type of OS_CANCEL : constant is 1;
end out_switch;
