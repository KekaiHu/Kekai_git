library verilog;
use verilog.vl_types.all;
entity DE4_Ethernet is
    port(
        GCLKIN          : in     vl_logic;
        GCLKOUT_FPGA    : out    vl_logic;
        OSC_50_BANK2    : in     vl_logic;
        OSC_50_BANK3    : in     vl_logic;
        OSC_50_BANK4    : in     vl_logic;
        OSC_50_BANK5    : in     vl_logic;
        OSC_50_BANK6    : in     vl_logic;
        OSC_50_BANK7    : in     vl_logic;
        PLL_CLKIN_p     : in     vl_logic;
        MAX_I2C_SCLK    : out    vl_logic;
        MAX_I2C_SDAT    : inout  vl_logic;
        LED             : out    vl_logic_vector(7 downto 0);
        BUTTON          : in     vl_logic_vector(3 downto 0);
        CPU_RESET_n     : in     vl_logic;
        EXT_IO          : inout  vl_logic;
        SW              : in     vl_logic_vector(7 downto 0);
        SLIDE_SW        : in     vl_logic_vector(3 downto 0);
        SEG0_D          : out    vl_logic_vector(6 downto 0);
        SEG0_DP         : out    vl_logic;
        SEG1_D          : out    vl_logic_vector(6 downto 0);
        SEG1_DP         : out    vl_logic;
        TEMP_INT_n      : in     vl_logic;
        TEMP_SMCLK      : out    vl_logic;
        TEMP_SMDAT      : inout  vl_logic;
        CSENSE_ADC_FO   : out    vl_logic;
        CSENSE_CS_n     : out    vl_logic_vector(1 downto 0);
        CSENSE_SCK      : out    vl_logic;
        CSENSE_SDI      : out    vl_logic;
        CSENSE_SDO      : in     vl_logic;
        FAN_CTRL        : out    vl_logic;
        EEP_SCL         : out    vl_logic;
        EEP_SDA         : inout  vl_logic;
        SD_CLK          : out    vl_logic;
        SD_CMD          : inout  vl_logic;
        SD_DAT          : inout  vl_logic_vector(3 downto 0);
        SD_WP_n         : in     vl_logic;
        UART_CTS        : out    vl_logic;
        UART_RTS        : in     vl_logic;
        UART_RXD        : in     vl_logic;
        UART_TXD        : out    vl_logic;
        ETH_INT_n       : in     vl_logic_vector(3 downto 0);
        ETH_MDC         : out    vl_logic_vector(3 downto 0);
        ETH_MDIO        : inout  vl_logic_vector(3 downto 0);
        ETH_RST_n       : out    vl_logic;
        ETH_RX_p        : in     vl_logic_vector(3 downto 0);
        ETH_TX_p        : out    vl_logic_vector(3 downto 0);
        PCIE_PREST_n    : in     vl_logic;
        PCIE_REFCLK_p   : in     vl_logic;
        PCIE_RX_p       : in     vl_logic;
        PCIE_SMBCLK     : in     vl_logic;
        PCIE_SMBDAT     : inout  vl_logic;
        PCIE_TX_p       : out    vl_logic;
        PCIE_WAKE_n     : out    vl_logic;
        FLASH_ADV_n     : out    vl_logic;
        FLASH_CLK       : out    vl_logic;
        FLASH_RESET_n   : out    vl_logic;
        FLASH_RYBY_n    : in     vl_logic;
        SSRAM_ADV       : out    vl_logic;
        SSRAM_BWA_n     : out    vl_logic;
        SSRAM_BWB_n     : out    vl_logic;
        SSRAM_CE_n      : out    vl_logic;
        SSRAM_CKE_n     : out    vl_logic;
        SSRAM_CLK       : out    vl_logic;
        SSRAM_OE_n      : out    vl_logic;
        SSRAM_WE_n      : out    vl_logic
    );
end DE4_Ethernet;
