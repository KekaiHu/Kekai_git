library verilog;
use verilog.vl_types.all;
entity output_queues is
    generic(
        DATA_WIDTH      : integer := 64;
        CTRL_WIDTH      : vl_notype;
        UDP_REG_SRC_WIDTH: integer := 2;
        OP_LUT_STAGE_NUM: integer := 4;
        NUM_OUTPUT_QUEUES: integer := 8;
        STAGE_NUM       : integer := 6;
        SRAM_ADDR_WIDTH : integer := 13
    );
    port(
        out_data_0      : out    vl_logic_vector;
        out_ctrl_0      : out    vl_logic_vector;
        out_rdy_0       : in     vl_logic;
        out_wr_0        : out    vl_logic;
        out_data_1      : out    vl_logic_vector;
        out_ctrl_1      : out    vl_logic_vector;
        out_rdy_1       : in     vl_logic;
        out_wr_1        : out    vl_logic;
        out_data_2      : out    vl_logic_vector;
        out_ctrl_2      : out    vl_logic_vector;
        out_rdy_2       : in     vl_logic;
        out_wr_2        : out    vl_logic;
        out_data_3      : out    vl_logic_vector;
        out_ctrl_3      : out    vl_logic_vector;
        out_rdy_3       : in     vl_logic;
        out_wr_3        : out    vl_logic;
        out_data_4      : out    vl_logic_vector;
        out_ctrl_4      : out    vl_logic_vector;
        out_rdy_4       : in     vl_logic;
        out_wr_4        : out    vl_logic;
        out_data_5      : out    vl_logic_vector;
        out_ctrl_5      : out    vl_logic_vector;
        out_wr_5        : out    vl_logic;
        out_rdy_5       : in     vl_logic;
        out_data_6      : out    vl_logic_vector;
        out_ctrl_6      : out    vl_logic_vector;
        out_wr_6        : out    vl_logic;
        out_rdy_6       : in     vl_logic;
        out_data_7      : out    vl_logic_vector;
        out_ctrl_7      : out    vl_logic_vector;
        out_wr_7        : out    vl_logic;
        out_rdy_7       : in     vl_logic;
        in_data         : in     vl_logic_vector;
        in_ctrl         : in     vl_logic_vector;
        in_rdy          : out    vl_logic;
        in_wr           : in     vl_logic;
        reg_req_in      : in     vl_logic;
        reg_ack_in      : in     vl_logic;
        reg_rd_wr_L_in  : in     vl_logic;
        reg_addr_in     : in     vl_logic_vector(22 downto 0);
        reg_data_in     : in     vl_logic_vector(31 downto 0);
        reg_src_in      : in     vl_logic_vector;
        reg_req_out     : out    vl_logic;
        reg_ack_out     : out    vl_logic;
        reg_rd_wr_L_out : out    vl_logic;
        reg_addr_out    : out    vl_logic_vector(22 downto 0);
        reg_data_out    : out    vl_logic_vector(31 downto 0);
        reg_src_out     : out    vl_logic_vector;
        wr_0_addr       : out    vl_logic_vector;
        wr_0_req        : out    vl_logic;
        wr_0_ack        : in     vl_logic;
        wr_0_data       : out    vl_logic_vector;
        rd_0_ack        : in     vl_logic;
        rd_0_data       : in     vl_logic_vector;
        rd_0_vld        : in     vl_logic;
        rd_0_addr       : out    vl_logic_vector;
        rd_0_req        : out    vl_logic;
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CTRL_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of UDP_REG_SRC_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of OP_LUT_STAGE_NUM : constant is 1;
    attribute mti_svvh_generic_type of NUM_OUTPUT_QUEUES : constant is 1;
    attribute mti_svvh_generic_type of STAGE_NUM : constant is 1;
    attribute mti_svvh_generic_type of SRAM_ADDR_WIDTH : constant is 1;
end output_queues;
