module state_machine(
input clk,
input [3:0] four_bit_hash,
input [11:0] pc_in,
input new_inst_signal,
input reset,
output packet_drop_signal
);


reg [10:0] state_reg,next_state;
wire [9:0] pc;
reg packet_drop_signal_register,packet_drop_signal_out;
	//`define 1000 = 1000;

	always @(posedge clk) begin	
		if (reset) begin
			state_reg <= 0; // initialize state reg to idle
			packet_drop_signal_out = 0;
		end
		else begin
			if(new_inst_signal)begin
				state_reg <= next_state;	
				packet_drop_signal_out = packet_drop_signal_register;
			end
		end
	end 
assign pc = pc_in[11:2];
	always@(*)begin

case(state_reg) 
//1999:begin if(four_bit_hash == 3) begin next_state = 0; end else begin next_state = 2000; end end
0: begin if(four_bit_hash == 0) next_state = 1; else  next_state = 2000;  end 
1: begin if(four_bit_hash == 7) next_state = 4; else if (four_bit_hash == 3) next_state = 2; else next_state = 2000;  end 
2: begin if(four_bit_hash == 0) next_state = 3; else  next_state = 2000;  end 
3: begin if(four_bit_hash == 4) next_state = 21; else if (four_bit_hash == 7) next_state = 4; else next_state = 2000;  end 
4: begin if(four_bit_hash == 11) next_state = 5; else  next_state = 2000;  end 
5: begin if(four_bit_hash == 5) next_state = 6; else  next_state = 2000;  end 
6: begin if(four_bit_hash == 7) next_state = 7; else  next_state = 2000;  end 
7: begin if(four_bit_hash == 6) next_state = 8; else  next_state = 2000;  end 
8: begin if(four_bit_hash == 10) next_state = 9; else  next_state = 2000;  end 
9: begin if(four_bit_hash == 8) next_state = 10; else  next_state = 2000;  end 
10: begin if(four_bit_hash == 5) next_state = 11; else  next_state = 2000;  end 
11: begin if(four_bit_hash == 5) next_state = 12; else  next_state = 2000;  end 
12: begin if(four_bit_hash == 8) next_state = 13; else  next_state = 2000;  end 
13: begin if(four_bit_hash == 3) next_state = 14; else  next_state = 2000;  end 
14: begin if(four_bit_hash == 5) next_state = 15; else  next_state = 2000;  end 
15: begin if(four_bit_hash == 5 && pc == 10'hc) next_state = 12; else if (four_bit_hash == 5 && pc == 10'h10) next_state = 16; else next_state = 2000;  end 
16: begin if(four_bit_hash == 5) next_state = 17; else  next_state = 2000;  end 
17: begin if(four_bit_hash == 6) next_state = 18; else  next_state = 2000;  end 
18: begin if(four_bit_hash == 0) next_state = 19; else  next_state = 2000;  end 
19: begin if(four_bit_hash == 5) next_state = 89; else if (four_bit_hash == 3) next_state = 20; else next_state = 2000;  end 
20: begin if(four_bit_hash == 4) next_state = 21; else  next_state = 2000;  end 
21: begin if(four_bit_hash == 3) next_state = 20; else if (four_bit_hash == 9) next_state = 22; else next_state = 2000;  end 
22: begin if(four_bit_hash == 10) next_state = 23; else  next_state = 2000;  end 
23: begin if(four_bit_hash == 11) next_state = 24; else  next_state = 2000;  end 
24: begin if(four_bit_hash == 11) next_state = 25; else  next_state = 2000;  end 
25: begin if(four_bit_hash == 12) next_state = 26; else  next_state = 2000;  end 
26: begin if(four_bit_hash == 13) next_state = 27; else  next_state = 2000;  end 
27: begin if(four_bit_hash == 12) next_state = 28; else  next_state = 2000;  end 
28: begin if(four_bit_hash == 11) next_state = 29; else  next_state = 2000;  end 
29: begin if(four_bit_hash == 12) next_state = 30; else  next_state = 2000;  end 
30: begin if(four_bit_hash == 13) next_state = 31; else  next_state = 2000;  end 
31: begin if(four_bit_hash == 13) next_state = 32; else  next_state = 2000;  end 
32: begin if(four_bit_hash == 13) next_state = 33; else  next_state = 2000;  end 
33: begin if(four_bit_hash == 15) next_state = 34; else  next_state = 2000;  end 
34: begin if(four_bit_hash == 15) next_state = 35; else  next_state = 2000;  end 
35: begin if(four_bit_hash == 13) next_state = 36; else  next_state = 2000;  end 
36: begin if(four_bit_hash == 11) next_state = 37; else  next_state = 2000;  end 
37: begin if(four_bit_hash == 12) next_state = 38; else  next_state = 2000;  end 
38: begin if(four_bit_hash == 13) next_state = 39; else  next_state = 2000;  end 
39: begin if(four_bit_hash == 13) next_state = 40; else  next_state = 2000;  end 
40: begin if(four_bit_hash == 13) next_state = 41; else  next_state = 2000;  end 
41: begin if(four_bit_hash == 14) next_state = 42; else  next_state = 2000;  end 
42: begin if(four_bit_hash == 15) next_state = 43; else  next_state = 2000;  end 
43: begin if(four_bit_hash == 14) next_state = 44; else  next_state = 2000;  end 
44: begin if(four_bit_hash == 13) next_state = 45; else  next_state = 2000;  end 
45: begin if(four_bit_hash == 14) next_state = 46; else  next_state = 2000;  end 
46: begin if(four_bit_hash == 1) next_state = 47; else  next_state = 2000;  end 
47: begin if(four_bit_hash == 5) next_state = 48; else  next_state = 2000;  end 
48: begin if(four_bit_hash == 0) next_state = 49; else  next_state = 2000;  end 
49: begin if(four_bit_hash == 7) next_state = 81; else if (four_bit_hash == 8) next_state = 50; else next_state = 2000;  end 
50: begin if(four_bit_hash == 9) next_state = 51; else  next_state = 2000;  end 
51: begin if(four_bit_hash == 10) next_state = 52; else  next_state = 2000;  end 
52: begin if(four_bit_hash == 10) next_state = 53; else  next_state = 2000;  end 
53: begin if(four_bit_hash == 11) next_state = 54; else  next_state = 2000;  end 
54: begin if(four_bit_hash == 12) next_state = 55; else  next_state = 2000;  end 
55: begin if(four_bit_hash == 11) next_state = 56; else  next_state = 2000;  end 
56: begin if(four_bit_hash == 10) next_state = 57; else  next_state = 2000;  end 
57: begin if(four_bit_hash == 11) next_state = 58; else  next_state = 2000;  end 
58: begin if(four_bit_hash == 12) next_state = 59; else  next_state = 2000;  end 
59: begin if(four_bit_hash == 12) next_state = 60; else  next_state = 2000;  end 
60: begin if(four_bit_hash == 12) next_state = 61; else  next_state = 2000;  end 
61: begin if(four_bit_hash == 14) next_state = 62; else  next_state = 2000;  end 
62: begin if(four_bit_hash == 14) next_state = 63; else  next_state = 2000;  end 
63: begin if(four_bit_hash == 12) next_state = 64; else  next_state = 2000;  end 
64: begin if(four_bit_hash == 10) next_state = 65; else  next_state = 2000;  end 
65: begin if(four_bit_hash == 11) next_state = 66; else  next_state = 2000;  end 
66: begin if(four_bit_hash == 12) next_state = 67; else  next_state = 2000;  end 
67: begin if(four_bit_hash == 12) next_state = 68; else  next_state = 2000;  end 
68: begin if(four_bit_hash == 12) next_state = 69; else  next_state = 2000;  end 
69: begin if(four_bit_hash == 13) next_state = 70; else  next_state = 2000;  end 
70: begin if(four_bit_hash == 14) next_state = 71; else  next_state = 2000;  end 
71: begin if(four_bit_hash == 13) next_state = 72; else  next_state = 2000;  end 
72: begin if(four_bit_hash == 12) next_state = 73; else  next_state = 2000;  end 
73: begin if(four_bit_hash == 13) next_state = 74; else  next_state = 2000;  end 
74: begin if(four_bit_hash == 0) next_state = 75; else  next_state = 2000;  end 
75: begin if(four_bit_hash == 13) next_state = 76; else  next_state = 2000;  end 
76: begin if(four_bit_hash == 7) next_state = 77; else  next_state = 2000;  end 
77: begin if(four_bit_hash == 8) next_state = 78; else  next_state = 2000;  end 
78: begin if(four_bit_hash == 5) next_state = 79; else  next_state = 2000;  end 
79: begin if(four_bit_hash == 7) next_state = 80; else  next_state = 2000;  end 
80: begin if(four_bit_hash == 7) next_state = 81; else  next_state = 2000;  end 
81: begin if(four_bit_hash == 13) next_state = 82; else  next_state = 2000;  end 
82: begin if(four_bit_hash == 10) next_state = 83; else  next_state = 2000;  end 
83: begin if(four_bit_hash == 10) next_state = 84; else  next_state = 2000;  end 
84: begin if(four_bit_hash == 12) next_state = 85; else  next_state = 2000;  end 
85: begin if(four_bit_hash == 11) next_state = 86; else  next_state = 2000;  end 
86: begin if(four_bit_hash == 6) next_state = 87; else  next_state = 2000;  end 
87: begin if(four_bit_hash == 0) next_state = 88; else  next_state = 2000;  end 
88: begin if(four_bit_hash == 5) next_state = 89; else  next_state = 2000;  end 
89: begin if(four_bit_hash == 15) next_state = 90; else  next_state = 2000;  end 
90: begin if(four_bit_hash == 10) next_state = 91; else  next_state = 2000;  end 
91: begin if(four_bit_hash == 12) next_state = 92; else  next_state = 2000;  end 
92: begin if(four_bit_hash == 14) next_state = 93; else  next_state = 2000;  end 
93: begin if(four_bit_hash == 9) next_state = 94; else  next_state = 2000;  end 
94: begin if(four_bit_hash == 14) next_state = 95; else  next_state = 2000;  end 
95: begin if(four_bit_hash == 9) next_state = 96; else  next_state = 2000;  end 
96: begin if(four_bit_hash == 9) next_state = 97; else  next_state = 2000;  end 
97: begin if(four_bit_hash == 7) next_state = 98; else  next_state = 2000;  end 
98: begin if(four_bit_hash == 6) next_state = 99; else  next_state = 2000;  end 
99: begin if(four_bit_hash == 7) next_state = 100; else  next_state = 2000;  end 
100: begin if(four_bit_hash == 5) next_state = 101; else  next_state = 2000;  end 
101: begin if(four_bit_hash == 0) next_state = 102; else  next_state = 2000;  end 
102: begin if(four_bit_hash == 8) next_state = 103; else  next_state = 2000;  end 
103: begin if(four_bit_hash == 7) next_state = 104; else  next_state = 2000;  end 
104: begin if(four_bit_hash == 0) next_state = 105; else  next_state = 2000;  end 
105: begin if(four_bit_hash == 4) next_state = 106; else  next_state = 2000;  end 
106: begin if(four_bit_hash == 11) next_state = 107; else  next_state = 2000;  end 
107: begin if(four_bit_hash == 11) next_state = 108; else  next_state = 2000;  end 
108: begin if(four_bit_hash == 4) next_state = 109; else  next_state = 2000;  end 
109: begin if(four_bit_hash == 11) next_state = 110; else  next_state = 2000;  end 
110: begin if(four_bit_hash == 0) next_state = 111; else  next_state = 2000;  end 
111: begin if(four_bit_hash == 13) next_state = 318; else if (four_bit_hash == 9) next_state = 112; else next_state = 2000;  end 
112: begin if(four_bit_hash == 6) next_state = 113; else  next_state = 2000;  end 
113: begin if(four_bit_hash == 8) next_state = 114; else  next_state = 2000;  end 
114: begin if(four_bit_hash == 5) next_state = 115; else  next_state = 2000;  end 
115: begin if(four_bit_hash == 0) next_state = 116; else  next_state = 2000;  end 
116: begin if(four_bit_hash == 8) next_state = 117; else  next_state = 2000;  end 
117: begin if(four_bit_hash == 7) next_state = 118; else  next_state = 2000;  end 
118: begin if(four_bit_hash == 0) next_state = 119; else  next_state = 2000;  end 
119: begin if(four_bit_hash == 12) next_state = 120; else  next_state = 2000;  end 
120: begin if(four_bit_hash == 4) next_state = 121; else  next_state = 2000;  end 
121: begin if(four_bit_hash == 10) next_state = 122; else  next_state = 2000;  end 
122: begin if(four_bit_hash == 9) next_state = 123; else  next_state = 2000;  end 
123: begin if(four_bit_hash == 0) next_state = 124; else  next_state = 2000;  end 
124: begin if(four_bit_hash == 4) next_state = 125; else  next_state = 2000;  end 
125: begin if(four_bit_hash == 0) next_state = 126; else  next_state = 2000;  end 
126: begin if(four_bit_hash == 13) next_state = 318; else if (four_bit_hash == 6) next_state = 127; else next_state = 2000;  end 
127: begin if(four_bit_hash == 7) next_state = 128; else  next_state = 2000;  end 
128: begin if(four_bit_hash == 5) next_state = 129; else  next_state = 2000;  end 
129: begin if(four_bit_hash == 0) next_state = 130; else  next_state = 2000;  end 
130: begin if(four_bit_hash == 8) next_state = 131; else  next_state = 2000;  end 
131: begin if(four_bit_hash == 7) next_state = 132; else  next_state = 2000;  end 
132: begin if(four_bit_hash == 0) next_state = 133; else  next_state = 2000;  end 
133: begin if(four_bit_hash == 4) next_state = 134; else  next_state = 2000;  end 
134: begin if(four_bit_hash == 12) next_state = 135; else  next_state = 2000;  end 
135: begin if(four_bit_hash == 6) next_state = 136; else  next_state = 2000;  end 
136: begin if(four_bit_hash == 7) next_state = 137; else  next_state = 2000;  end 
137: begin if(four_bit_hash == 5) next_state = 138; else  next_state = 2000;  end 
138: begin if(four_bit_hash == 0) next_state = 139; else  next_state = 2000;  end 
139: begin if(four_bit_hash == 8) next_state = 140; else  next_state = 2000;  end 
140: begin if(four_bit_hash == 7) next_state = 141; else  next_state = 2000;  end 
141: begin if(four_bit_hash == 0) next_state = 142; else  next_state = 2000;  end 
142: begin if(four_bit_hash == 4) next_state = 143; else  next_state = 2000;  end 
143: begin if(four_bit_hash == 12) next_state = 144; else  next_state = 2000;  end 
144: begin if(four_bit_hash == 11) next_state = 145; else  next_state = 2000;  end 
145: begin if(four_bit_hash == 0) next_state = 146; else  next_state = 2000;  end 
146: begin if(four_bit_hash == 3) next_state = 147; else  next_state = 2000;  end 
147: begin if(four_bit_hash == 10) next_state = 148; else  next_state = 2000;  end 
148: begin if(four_bit_hash == 10) next_state = 149; else  next_state = 2000;  end 
149: begin if(four_bit_hash == 11) next_state = 150; else  next_state = 2000;  end 
150: begin if(four_bit_hash == 0) next_state = 151; else  next_state = 2000;  end 
151: begin if(four_bit_hash == 6) next_state = 152; else  next_state = 2000;  end 
152: begin if(four_bit_hash == 11) next_state = 153; else  next_state = 2000;  end 
153: begin if(four_bit_hash == 10) next_state = 154; else  next_state = 2000;  end 
154: begin if(four_bit_hash == 13) next_state = 155; else  next_state = 2000;  end 
155: begin if(four_bit_hash == 7) next_state = 156; else  next_state = 2000;  end 
156: begin if(four_bit_hash == 10) next_state = 157; else  next_state = 2000;  end 
157: begin if(four_bit_hash == 0) next_state = 158; else  next_state = 2000;  end 
158: begin if(four_bit_hash == 7) next_state = 159; else  next_state = 2000;  end 
159: begin if(four_bit_hash == 9) next_state = 160; else  next_state = 2000;  end 
160: begin if(four_bit_hash == 6) next_state = 161; else  next_state = 2000;  end 
161: begin if(four_bit_hash == 0) next_state = 162; else  next_state = 2000;  end 
162: begin if(four_bit_hash == 9) next_state = 220; else if (four_bit_hash == 13) next_state = 163; else next_state = 2000;  end 
163: begin if(four_bit_hash == 8) next_state = 164; else  next_state = 2000;  end 
164: begin if(four_bit_hash == 10) next_state = 165; else  next_state = 2000;  end 
165: begin if(four_bit_hash == 0) next_state = 166; else  next_state = 2000;  end 
166: begin if(four_bit_hash == 7) next_state = 167; else  next_state = 2000;  end 
167: begin if(four_bit_hash == 10) next_state = 168; else  next_state = 2000;  end 
168: begin if(four_bit_hash == 9) next_state = 169; else  next_state = 2000;  end 
169: begin if(four_bit_hash == 9) next_state = 170; else  next_state = 2000;  end 
170: begin if(four_bit_hash == 6) next_state = 171; else  next_state = 2000;  end 
171: begin if(four_bit_hash == 3) next_state = 172; else  next_state = 2000;  end 
172: begin if(four_bit_hash == 10) next_state = 173; else  next_state = 2000;  end 
173: begin if(four_bit_hash == 5) next_state = 174; else  next_state = 2000;  end 
174: begin if(four_bit_hash == 5) next_state = 175; else  next_state = 2000;  end 
175: begin if(four_bit_hash == 0) next_state = 176; else  next_state = 2000;  end 
176: begin if(four_bit_hash == 12) next_state = 177; else  next_state = 2000;  end 
177: begin if(four_bit_hash == 10) next_state = 178; else  next_state = 2000;  end 
178: begin if(four_bit_hash == 9) next_state = 179; else  next_state = 2000;  end 
179: begin if(four_bit_hash == 6) next_state = 180; else  next_state = 2000;  end 
180: begin if(four_bit_hash == 3) next_state = 181; else  next_state = 2000;  end 
181: begin if(four_bit_hash == 10) next_state = 182; else  next_state = 2000;  end 
182: begin if(four_bit_hash == 5) next_state = 183; else  next_state = 2000;  end 
183: begin if(four_bit_hash == 5) next_state = 184; else  next_state = 2000;  end 
184: begin if(four_bit_hash == 0) next_state = 185; else  next_state = 2000;  end 
185: begin if(four_bit_hash == 4) next_state = 186; else  next_state = 2000;  end 
186: begin if(four_bit_hash == 11) next_state = 187; else  next_state = 2000;  end 
187: begin if(four_bit_hash == 10) next_state = 188; else  next_state = 2000;  end 
188: begin if(four_bit_hash == 0) next_state = 189; else  next_state = 2000;  end 
189: begin if(four_bit_hash == 5) next_state = 190; else  next_state = 2000;  end 
190: begin if(four_bit_hash == 10) next_state = 191; else  next_state = 2000;  end 
191: begin if(four_bit_hash == 0) next_state = 192; else  next_state = 2000;  end 
192: begin if(four_bit_hash == 8) next_state = 193; else  next_state = 2000;  end 
193: begin if(four_bit_hash == 0) next_state = 194; else  next_state = 2000;  end 
194: begin if(four_bit_hash == 9) next_state = 216; else if (four_bit_hash == 4) next_state = 195; else next_state = 2000;  end 
195: begin if(four_bit_hash == 11) next_state = 196; else  next_state = 2000;  end 
196: begin if(four_bit_hash == 9) next_state = 197; else  next_state = 2000;  end 
197: begin if(four_bit_hash == 0) next_state = 198; else  next_state = 2000;  end 
198: begin if(four_bit_hash == 3) next_state = 199; else  next_state = 2000;  end 
199: begin if(four_bit_hash == 10) next_state = 200; else  next_state = 2000;  end 
200: begin if(four_bit_hash == 6) next_state = 201; else  next_state = 2000;  end 
201: begin if(four_bit_hash == 5) next_state = 202; else  next_state = 2000;  end 
202: begin if(four_bit_hash == 0) next_state = 203; else  next_state = 2000;  end 
203: begin if(four_bit_hash == 11) next_state = 204; else  next_state = 2000;  end 
204: begin if(four_bit_hash == 11) next_state = 205; else  next_state = 2000;  end 
205: begin if(four_bit_hash == 9) next_state = 206; else  next_state = 2000;  end 
206: begin if(four_bit_hash == 0) next_state = 207; else  next_state = 2000;  end 
207: begin if(four_bit_hash == 7) next_state = 208; else  next_state = 2000;  end 
208: begin if(four_bit_hash == 11) next_state = 209; else  next_state = 2000;  end 
209: begin if(four_bit_hash == 7) next_state = 210; else  next_state = 2000;  end 
210: begin if(four_bit_hash == 10) next_state = 211; else  next_state = 2000;  end 
211: begin if(four_bit_hash == 0) next_state = 212; else  next_state = 2000;  end 
212: begin if(four_bit_hash == 7) next_state = 213; else  next_state = 2000;  end 
213: begin if(four_bit_hash == 5) next_state = 214; else  next_state = 2000;  end 
214: begin if(four_bit_hash == 0) next_state = 215; else  next_state = 2000;  end 
215: begin if(four_bit_hash == 13) next_state = 225; else if (four_bit_hash == 9) next_state = 216; else next_state = 2000;  end 
216: begin if(four_bit_hash == 0) next_state = 217; else  next_state = 2000;  end 
217: begin if(four_bit_hash == 5) next_state = 218; else  next_state = 2000;  end 
218: begin if(four_bit_hash == 10) next_state = 219; else  next_state = 2000;  end 
219: begin if(four_bit_hash == 9) next_state = 220; else  next_state = 2000;  end 
220: begin if(four_bit_hash == 0) next_state = 221; else  next_state = 2000;  end 
221: begin if(four_bit_hash == 8) next_state = 222; else  next_state = 2000;  end 
222: begin if(four_bit_hash == 15) next_state = 223; else  next_state = 2000;  end 
223: begin if(four_bit_hash == 0) next_state = 224; else  next_state = 2000;  end 
224: begin if(four_bit_hash == 13 && pc == 163) next_state = 163; else if (four_bit_hash == 13 && pc == 225) next_state = 225; else next_state = 2000;  end 
225: begin if(four_bit_hash == 7) next_state = 226; else  next_state = 2000;  end 
226: begin if(four_bit_hash == 9) next_state = 227; else  next_state = 2000;  end 
227: begin if(four_bit_hash == 0) next_state = 228; else  next_state = 2000;  end 
228: begin if(four_bit_hash == 7) next_state = 229; else  next_state = 2000;  end 
229: begin if(four_bit_hash == 10) next_state = 230; else  next_state = 2000;  end 
230: begin if(four_bit_hash == 0) next_state = 231; else  next_state = 2000;  end 
231: begin if(four_bit_hash == 6) next_state = 232; else  next_state = 2000;  end 
232: begin if(four_bit_hash == 0) next_state = 233; else  next_state = 2000;  end 
233: begin if(four_bit_hash == 9) next_state = 246; else if (four_bit_hash == 6) next_state = 234; else next_state = 2000;  end 
234: begin if(four_bit_hash == 5) next_state = 235; else  next_state = 2000;  end 
235: begin if(four_bit_hash == 0) next_state = 236; else  next_state = 2000;  end 
236: begin if(four_bit_hash == 11) next_state = 237; else  next_state = 2000;  end 
237: begin if(four_bit_hash == 11) next_state = 238; else  next_state = 2000;  end 
238: begin if(four_bit_hash == 6) next_state = 239; else  next_state = 2000;  end 
239: begin if(four_bit_hash == 7) next_state = 240; else  next_state = 2000;  end 
240: begin if(four_bit_hash == 11) next_state = 241; else  next_state = 2000;  end 
241: begin if(four_bit_hash == 7) next_state = 242; else  next_state = 2000;  end 
242: begin if(four_bit_hash == 10) next_state = 243; else  next_state = 2000;  end 
243: begin if(four_bit_hash == 0) next_state = 244; else  next_state = 2000;  end 
244: begin if(four_bit_hash == 7) next_state = 245; else  next_state = 2000;  end 
245: begin if(four_bit_hash == 9) next_state = 246; else  next_state = 2000;  end 
246: begin if(four_bit_hash == 0) next_state = 247; else  next_state = 2000;  end 
247: begin if(four_bit_hash == 4) next_state = 248; else  next_state = 2000;  end 
248: begin if(four_bit_hash == 10) next_state = 249; else  next_state = 2000;  end 
249: begin if(four_bit_hash == 6) next_state = 250; else  next_state = 2000;  end 
250: begin if(four_bit_hash == 8) next_state = 251; else  next_state = 2000;  end 
251: begin if(four_bit_hash == 5) next_state = 252; else  next_state = 2000;  end 
252: begin if(four_bit_hash == 0) next_state = 253; else  next_state = 2000;  end 
253: begin if(four_bit_hash == 8) next_state = 254; else  next_state = 2000;  end 
254: begin if(four_bit_hash == 8) next_state = 255; else  next_state = 2000;  end 
255: begin if(four_bit_hash == 5) next_state = 256; else  next_state = 2000;  end 
256: begin if(four_bit_hash == 13) next_state = 257; else  next_state = 2000;  end 
257: begin if(four_bit_hash == 6) next_state = 258; else  next_state = 2000;  end 
258: begin if(four_bit_hash == 8) next_state = 259; else  next_state = 2000;  end 
259: begin if(four_bit_hash == 9) next_state = 260; else  next_state = 2000;  end 
260: begin if(four_bit_hash == 0) next_state = 261; else  next_state = 2000;  end 
261: begin if(four_bit_hash == 4) next_state = 262; else  next_state = 2000;  end 
262: begin if(four_bit_hash == 7) next_state = 263; else  next_state = 2000;  end 
263: begin if(four_bit_hash == 0) next_state = 264; else  next_state = 2000;  end 
264: begin if(four_bit_hash == 7) next_state = 265; else  next_state = 2000;  end 
265: begin if(four_bit_hash == 8) next_state = 266; else  next_state = 2000;  end 
266: begin if(four_bit_hash == 6) next_state = 267; else  next_state = 2000;  end 
267: begin if(four_bit_hash == 9) next_state = 268; else  next_state = 2000;  end 
268: begin if(four_bit_hash == 7) next_state = 269; else  next_state = 2000;  end 
269: begin if(four_bit_hash == 0) next_state = 270; else  next_state = 2000;  end 
270: begin if(four_bit_hash == 7) next_state = 271; else  next_state = 2000;  end 
271: begin if(four_bit_hash == 8) next_state = 272; else  next_state = 2000;  end 
272: begin if(four_bit_hash == 6) next_state = 273; else  next_state = 2000;  end 
273: begin if(four_bit_hash == 6) next_state = 274; else  next_state = 2000;  end 
274: begin if(four_bit_hash == 5) next_state = 275; else  next_state = 2000;  end 
275: begin if(four_bit_hash == 0) next_state = 276; else  next_state = 2000;  end 
276: begin if(four_bit_hash == 8) next_state = 277; else  next_state = 2000;  end 
277: begin if(four_bit_hash == 7) next_state = 278; else  next_state = 2000;  end 
278: begin if(four_bit_hash == 0) next_state = 279; else  next_state = 2000;  end 
279: begin if(four_bit_hash == 4) next_state = 280; else  next_state = 2000;  end 
280: begin if(four_bit_hash == 9) next_state = 281; else  next_state = 2000;  end 
281: begin if(four_bit_hash == 9) next_state = 282; else  next_state = 2000;  end 
282: begin if(four_bit_hash == 3) next_state = 283; else  next_state = 2000;  end 
283: begin if(four_bit_hash == 8) next_state = 284; else  next_state = 2000;  end 
284: begin if(four_bit_hash == 6) next_state = 285; else  next_state = 2000;  end 
285: begin if(four_bit_hash == 0) next_state = 286; else  next_state = 2000;  end 
286: begin if(four_bit_hash == 8 && pc == 293) next_state = 293; else if (four_bit_hash == 8 && pc == 287) next_state = 287; else next_state = 2000;  end 
287: begin if(four_bit_hash == 0) next_state = 288; else  next_state = 2000;  end 
288: begin if(four_bit_hash == 6) next_state = 289; else  next_state = 2000;  end 
289: begin if(four_bit_hash == 9) next_state = 290; else  next_state = 2000;  end 
290: begin if(four_bit_hash == 5) next_state = 291; else  next_state = 2000;  end 
291: begin if(four_bit_hash == 0) next_state = 292; else  next_state = 2000;  end 
292: begin if(four_bit_hash == 6) next_state = 297; else if (four_bit_hash == 8) next_state = 293; else next_state = 2000;  end 
293: begin if(four_bit_hash == 0) next_state = 294; else  next_state = 2000;  end 
294: begin if(four_bit_hash == 5) next_state = 295; else  next_state = 2000;  end 
295: begin if(four_bit_hash == 9) next_state = 296; else  next_state = 2000;  end 
296: begin if(four_bit_hash == 6) next_state = 297; else  next_state = 2000;  end 
297: begin if(four_bit_hash == 6) next_state = 298; else  next_state = 2000;  end 
298: begin if(four_bit_hash == 5) next_state = 299; else  next_state = 2000;  end 
299: begin if(four_bit_hash == 0) next_state = 300; else  next_state = 2000;  end 
300: begin if(four_bit_hash == 8) next_state = 301; else  next_state = 2000;  end 
301: begin if(four_bit_hash == 7) next_state = 302; else  next_state = 2000;  end 
302: begin if(four_bit_hash == 0) next_state = 303; else  next_state = 2000;  end 
303: begin if(four_bit_hash == 4) next_state = 304; else  next_state = 2000;  end 
304: begin if(four_bit_hash == 8) next_state = 305; else  next_state = 2000;  end 
305: begin if(four_bit_hash == 8) next_state = 306; else  next_state = 2000;  end 
306: begin if(four_bit_hash == 0) next_state = 307; else  next_state = 2000;  end 
307: begin if(four_bit_hash == 4) next_state = 308; else  next_state = 2000;  end 
308: begin if(four_bit_hash == 7) next_state = 309; else  next_state = 2000;  end 
309: begin if(four_bit_hash == 0) next_state = 310; else  next_state = 2000;  end 
310: begin if(four_bit_hash == 7) next_state = 311; else  next_state = 2000;  end 
311: begin if(four_bit_hash == 8) next_state = 312; else  next_state = 2000;  end 
312: begin if(four_bit_hash == 6) next_state = 313; else  next_state = 2000;  end 
313: begin if(four_bit_hash == 7) next_state = 314; else  next_state = 2000;  end 
314: begin if(four_bit_hash == 7) next_state = 315; else  next_state = 2000;  end 
315: begin if(four_bit_hash == 0) next_state = 316; else  next_state = 2000;  end 
316: begin if(four_bit_hash == 7) next_state = 317; else  next_state = 2000;  end 
317: begin if(four_bit_hash == 13) next_state = 318; else  next_state = 2000;  end 
318: begin if(four_bit_hash == 8) next_state = 319; else  next_state = 2000;  end 
319: begin if(four_bit_hash == 9) next_state = 320; else  next_state = 2000;  end 
320: begin if(four_bit_hash == 0) next_state = 321; else  next_state = 2000;  end 
321: begin if(four_bit_hash == 7) next_state = 322; else  next_state = 2000;  end 
322: begin if(four_bit_hash == 7) next_state = 323; else  next_state = 2000;  end 
323: begin if(four_bit_hash == 4) next_state = 324; else  next_state = 2000;  end 
324: begin if(four_bit_hash == 7) next_state = 325; else  next_state = 2000;  end 
325: begin if(four_bit_hash == 7) next_state = 326; else  next_state = 2000;  end 
326: begin if(four_bit_hash == 0) next_state = 327; else  next_state = 2000;  end 
327: begin if(four_bit_hash == 14) next_state = 95; else if (four_bit_hash == 0) next_state = 328; else next_state = 2000;  end 
328: begin if(four_bit_hash == 0) next_state = 329; else  next_state = 2000;  end 
329: begin if(four_bit_hash == 0) next_state = 330; else  next_state = 2000;  end 
330: begin if(four_bit_hash == 0) next_state = 331; else  next_state = 2000;  end 
331: begin if(four_bit_hash == 0) next_state = 332; else  next_state = 2000;  end 
332: begin if(four_bit_hash == 0) next_state = 333; else  next_state = 2000;  end 
333: begin if(four_bit_hash == 0) next_state = 334; else  next_state = 2000;  end 
334: begin if(four_bit_hash == 0) next_state = 335; else  next_state = 2000;  end 
335: begin if(four_bit_hash == 0) next_state = 336; else  next_state = 2000;  end 
336: begin if(four_bit_hash == 0) next_state = 337; else  next_state = 2000;  end 
337: begin if(four_bit_hash == 0) next_state = 338; else  next_state = 2000;  end 
338: begin if(four_bit_hash == 0) next_state = 339; else  next_state = 2000;  end 
339: begin if(four_bit_hash == 0) next_state = 340; else  next_state = 2000;  end 
340: begin if(four_bit_hash == 0) next_state = 341; else  next_state = 2000;  end 
341: begin if(four_bit_hash == 0) next_state = 342; else  next_state = 2000;  end 
342: begin if(four_bit_hash == 0) next_state = 343; else  next_state = 2000;  end 
343: begin if(four_bit_hash == 0) next_state = 344; else  next_state = 2000;  end 
344: begin if(four_bit_hash == 0) next_state = 345; else  next_state = 2000;  end 
345: begin if(four_bit_hash == 0) next_state = 346; else  next_state = 2000;  end 
346: begin if(four_bit_hash == 0) next_state = 347; else  next_state = 2000;  end 
347: begin if(four_bit_hash == 0) next_state = 348; else  next_state = 2000;  end 
348: begin if(four_bit_hash == 0) next_state = 349; else  next_state = 2000;  end 
349: begin if(four_bit_hash == 0) next_state = 350; else  next_state = 2000;  end 
350: begin if(four_bit_hash == 0) next_state = 351; else  next_state = 2000;  end 
351: begin if(four_bit_hash == 0) next_state = 352; else  next_state = 2000;  end 
352: begin if(four_bit_hash == 0) next_state = 353; else  next_state = 2000;  end 
353: begin if(four_bit_hash == 0) next_state = 354; else  next_state = 2000;  end 
354: begin if(four_bit_hash == 0) next_state = 355; else  next_state = 2000;  end 
355: begin if(four_bit_hash == 0) next_state = 356; else  next_state = 2000;  end 
356: begin if(four_bit_hash == 4) next_state = 357; else  next_state = 2000;  end 
357: begin if(four_bit_hash == 4) next_state = 358; else  next_state = 2000;  end 
358: begin if(four_bit_hash == 4) next_state = 359; else  next_state = 2000;  end 
359: begin if(four_bit_hash == 4) next_state = 360; else  next_state = 2000;  end 
360: begin if(four_bit_hash == 4) next_state = 361; else  next_state = 2000;  end 
361: begin if(four_bit_hash == 4) next_state = 362; else  next_state = 2000;  end 
362: begin if(four_bit_hash == 4) next_state = 363; else  next_state = 2000;  end 
363: begin if(four_bit_hash == 4) next_state = 364; else  next_state = 2000;  end 
364: begin if(four_bit_hash == 4) next_state = 365; else  next_state = 2000;  end 
365: begin if(four_bit_hash == 7) next_state = 366; else  next_state = 2000;  end 
366: begin if(four_bit_hash == 5) next_state = 367; else  next_state = 2000;  end 
367: begin if(four_bit_hash == 7) next_state = 368; else  next_state = 2000;  end 
368: begin if(four_bit_hash == 10) next_state = 369; else  next_state = 2000;  end 
369: begin if(four_bit_hash == 10) next_state = 370; else  next_state = 2000;  end 
370: begin if(four_bit_hash == 13) next_state = 371; else  next_state = 2000;  end 
371: begin if(four_bit_hash == 6) next_state = 372; else  next_state = 2000;  end 
372: begin if(four_bit_hash == 6) next_state = 373; else  next_state = 2000;  end 
373: begin if(four_bit_hash == 9) next_state = 374; else  next_state = 2000;  end 
374: begin if(four_bit_hash == 5) next_state = 375; else  next_state = 2000;  end 
375: begin if(four_bit_hash == 6) next_state = 376; else  next_state = 2000;  end 
376: begin if(four_bit_hash == 6) next_state = 377; else  next_state = 2000;  end 
377: begin if(four_bit_hash == 12) next_state = 378; else  next_state = 2000;  end 
378: begin if(four_bit_hash == 6) next_state = 379; else  next_state = 2000;  end 
379: begin if(four_bit_hash == 9) next_state = 380; else  next_state = 2000;  end 
380: begin if(four_bit_hash == 9) next_state = 381; else  next_state = 2000;  end 
381: begin if(four_bit_hash == 12) next_state = 382; else  next_state = 2000;  end 
382: begin if(four_bit_hash == 9) next_state = 383; else  next_state = 2000;  end 
383: begin if(four_bit_hash == 12) next_state = 384; else  next_state = 2000;  end 
384: begin if(four_bit_hash == 5) next_state = 385; else  next_state = 2000;  end 
385: begin if(four_bit_hash == 6) next_state = 386; else  next_state = 2000;  end 
386: begin if(four_bit_hash == 6) next_state = 387; else  next_state = 2000;  end 
387: begin if(four_bit_hash == 6) next_state = 388; else  next_state = 2000;  end 
388: begin if(four_bit_hash == 9) next_state = 389; else  next_state = 2000;  end 
389: begin if(four_bit_hash == 6) next_state = 390; else  next_state = 2000;  end 
390: begin if(four_bit_hash == 9) next_state = 391; else  next_state = 2000;  end 
391: begin if(four_bit_hash == 9) next_state = 392; else  next_state = 2000;  end 
392: begin if(four_bit_hash == 12) next_state = 393; else  next_state = 2000;  end 
393: begin if(four_bit_hash == 6) next_state = 394; else  next_state = 2000;  end 
394: begin if(four_bit_hash == 6) next_state = 395; else  next_state = 2000;  end 
395: begin if(four_bit_hash == 7) next_state = 396; else  next_state = 2000;  end 
396: begin if(four_bit_hash == 7) next_state = 397; else  next_state = 2000;  end 
397: begin if(four_bit_hash == 9) next_state = 398; else  next_state = 2000;  end 
398: begin if(four_bit_hash == 12) next_state = 399; else  next_state = 2000;  end 
399: begin if(four_bit_hash == 12) next_state = 400; else  next_state = 2000;  end 
400: begin if(four_bit_hash == 15) next_state = 401; else  next_state = 2000;  end 
401: begin if(four_bit_hash == 8) next_state = 402; else  next_state = 2000;  end 
402: begin if(four_bit_hash == 8) next_state = 403; else  next_state = 2000;  end 
403: begin if(four_bit_hash == 11) next_state = 404; else  next_state = 2000;  end 
404: begin if(four_bit_hash == 5) next_state = 405; else  next_state = 2000;  end 
405: begin if(four_bit_hash == 6) next_state = 406; else  next_state = 2000;  end 
406: begin if(four_bit_hash == 6) next_state = 407; else  next_state = 2000;  end 
407: begin if(four_bit_hash == 14) next_state = 408; else  next_state = 2000;  end 
408: begin if(four_bit_hash == 8) next_state = 409; else  next_state = 2000;  end 
409: begin if(four_bit_hash == 11) next_state = 410; else  next_state = 2000;  end 
410: begin if(four_bit_hash == 11) next_state = 411; else  next_state = 2000;  end 
411: begin if(four_bit_hash == 14) next_state = 412; else  next_state = 2000;  end 
412: begin if(four_bit_hash == 11) next_state = 413; else  next_state = 2000;  end 
413: begin if(four_bit_hash == 14) next_state = 414; else  next_state = 2000;  end 
414: begin if(four_bit_hash == 6) next_state = 415; else  next_state = 2000;  end 
415: begin if(four_bit_hash == 7) next_state = 416; else  next_state = 2000;  end 
416: begin if(four_bit_hash == 7) next_state = 417; else  next_state = 2000;  end 
417: begin if(four_bit_hash == 6) next_state = 418; else  next_state = 2000;  end 
418: begin if(four_bit_hash == 9) next_state = 419; else  next_state = 2000;  end 
419: begin if(four_bit_hash == 6) next_state = 420; else  next_state = 2000;  end 
420: begin if(four_bit_hash == 9) next_state = 421; else  next_state = 2000;  end 
421: begin if(four_bit_hash == 9) next_state = 422; else  next_state = 2000;  end 
422: begin if(four_bit_hash == 12) next_state = 423; else  next_state = 2000;  end 
423: begin if(four_bit_hash == 6) next_state = 424; else  next_state = 2000;  end 
424: begin if(four_bit_hash == 6) next_state = 425; else  next_state = 2000;  end 
425: begin if(four_bit_hash == 7) next_state = 426; else  next_state = 2000;  end 
426: begin if(four_bit_hash == 7) next_state = 427; else  next_state = 2000;  end 
427: begin if(four_bit_hash == 9) next_state = 428; else  next_state = 2000;  end 
428: begin if(four_bit_hash == 12) next_state = 429; else  next_state = 2000;  end 
429: begin if(four_bit_hash == 12) next_state = 430; else  next_state = 2000;  end 
430: begin if(four_bit_hash == 15) next_state = 431; else  next_state = 2000;  end 
431: begin if(four_bit_hash == 8) next_state = 432; else  next_state = 2000;  end 
432: begin if(four_bit_hash == 8) next_state = 433; else  next_state = 2000;  end 
433: begin if(four_bit_hash == 11) next_state = 434; else  next_state = 2000;  end 
434: begin if(four_bit_hash == 7) next_state = 435; else  next_state = 2000;  end 
435: begin if(four_bit_hash == 8) next_state = 436; else  next_state = 2000;  end 
436: begin if(four_bit_hash == 8) next_state = 437; else  next_state = 2000;  end 
437: begin if(four_bit_hash == 14) next_state = 438; else  next_state = 2000;  end 
438: begin if(four_bit_hash == 8) next_state = 439; else  next_state = 2000;  end 
439: begin if(four_bit_hash == 11) next_state = 440; else  next_state = 2000;  end 
440: begin if(four_bit_hash == 11) next_state = 441; else  next_state = 2000;  end 
441: begin if(four_bit_hash == 14) next_state = 442; else  next_state = 2000;  end 
442: begin if(four_bit_hash == 11) next_state = 443; else  next_state = 2000;  end 
443: begin if(four_bit_hash == 14) next_state = 444; else  next_state = 2000;  end 
444: begin if(four_bit_hash == 5) next_state = 445; else  next_state = 2000;  end 
445: begin if(four_bit_hash == 6) next_state = 446; else  next_state = 2000;  end 
446: begin if(four_bit_hash == 6) next_state = 447; else  next_state = 2000;  end 
447: begin if(four_bit_hash == 8) next_state = 448; else  next_state = 2000;  end 
448: begin if(four_bit_hash == 11) next_state = 449; else  next_state = 2000;  end 
449: begin if(four_bit_hash == 8) next_state = 450; else  next_state = 2000;  end 
450: begin if(four_bit_hash == 11) next_state = 451; else  next_state = 2000;  end 
451: begin if(four_bit_hash == 11) next_state = 452; else  next_state = 2000;  end 
452: begin if(four_bit_hash == 14) next_state = 453; else  next_state = 2000;  end 
453: begin if(four_bit_hash == 8) next_state = 454; else  next_state = 2000;  end 
454: begin if(four_bit_hash == 11) next_state = 455; else  next_state = 2000;  end 
455: begin if(four_bit_hash == 11) next_state = 456; else  next_state = 2000;  end 
456: begin if(four_bit_hash == 14) next_state = 457; else  next_state = 2000;  end 
457: begin if(four_bit_hash == 0) next_state = 458; else  next_state = 2000;  end 
458: begin if(four_bit_hash == 0) next_state = 459; else  next_state = 2000;  end 
459: begin if(four_bit_hash == 0) next_state = 460; else  next_state = 2000;  end 
460: begin if(four_bit_hash == 0) next_state = 461; else  next_state = 2000;  end 
461: begin if(four_bit_hash == 0) next_state = 462; else  next_state = 2000;  end 
462: begin if(four_bit_hash == 0) next_state = 463; else  next_state = 2000;  end 
463: begin if(four_bit_hash == 0) next_state = 464; else  next_state = 2000;  end 
464: begin if(four_bit_hash == 0) next_state = 465; else  next_state = 2000;  end 
465: begin if(four_bit_hash == 0) next_state = 466; else  next_state = 2000;  end 
466: begin if(four_bit_hash == 0) next_state = 467; else  next_state = 2000;  end 
467: begin if(four_bit_hash == 0) next_state = 468; else  next_state = 2000;  end 
468: begin if(four_bit_hash == 0) next_state = 469; else  next_state = 2000;  end 
469: begin if(four_bit_hash == 0) next_state = 470; else  next_state = 2000;  end 
470: begin if(four_bit_hash == 0) next_state = 471; else  next_state = 2000;  end 
471: begin if(four_bit_hash == 0) next_state = 472; else  next_state = 2000;  end 
472: begin if(four_bit_hash == 0) next_state = 473; else  next_state = 2000;  end 
473: begin if(four_bit_hash == 0) next_state = 474; else  next_state = 2000;  end 
474: begin if(four_bit_hash == 0) next_state = 475; else  next_state = 2000;  end 
475: begin if(four_bit_hash == 0) next_state = 476; else  next_state = 2000;  end 
476: begin if(four_bit_hash == 0) next_state = 477; else  next_state = 2000;  end 
477: begin if(four_bit_hash == 0) next_state = 478; else  next_state = 2000;  end 
478: begin if(four_bit_hash == 0) next_state = 479; else  next_state = 2000;  end 
479: begin if(four_bit_hash == 0) next_state = 480; else  next_state = 2000;  end 
480: begin if(four_bit_hash == 0) next_state = 481; else  next_state = 2000;  end 
481: begin if(four_bit_hash == 0) next_state = 482; else  next_state = 2000;  end 
482: begin if(four_bit_hash == 0) next_state = 483; else  next_state = 2000;  end 
483: begin if(four_bit_hash == 0) next_state = 484; else  next_state = 2000;  end 
484: begin if(four_bit_hash == 0) next_state = 485; else  next_state = 2000;  end 
485: begin if(four_bit_hash == 0) next_state = 486; else  next_state = 2000;  end 
486: begin if(four_bit_hash == 0) next_state = 487; else  next_state = 2000;  end 
487: begin if(four_bit_hash == 0) next_state = 488; else  next_state = 2000;  end 
488: begin if(four_bit_hash == 0) next_state = 489; else  next_state = 2000;  end 
489: begin if(four_bit_hash == 0) next_state = 490; else  next_state = 2000;  end 
490: begin if(four_bit_hash == 0) next_state = 491; else  next_state = 2000;  end 
491: begin if(four_bit_hash == 0) next_state = 492; else  next_state = 2000;  end 
492: begin if(four_bit_hash == 0) next_state = 493; else  next_state = 2000;  end 
493: begin if(four_bit_hash == 0) next_state = 494; else  next_state = 2000;  end 
494: begin if(four_bit_hash == 0) next_state = 495; else  next_state = 2000;  end 
495: begin if(four_bit_hash == 0) next_state = 496; else  next_state = 2000;  end 
496: begin if(four_bit_hash == 0) next_state = 497; else  next_state = 2000;  end 
497: begin if(four_bit_hash == 0) next_state = 498; else  next_state = 2000;  end 
498: begin if(four_bit_hash == 0) next_state = 499; else  next_state = 2000;  end 
499: begin if(four_bit_hash == 0) next_state = 500; else  next_state = 2000;  end 
500: begin if(four_bit_hash == 0) next_state = 501; else  next_state = 2000;  end 
501: begin if(four_bit_hash == 0) next_state = 502; else  next_state = 2000;  end 
502: begin if(four_bit_hash == 0) next_state = 503; else  next_state = 2000;  end 
503: begin if(four_bit_hash == 0) next_state = 504; else  next_state = 2000;  end 
504: begin if(four_bit_hash == 0) next_state = 505; else  next_state = 2000;  end 
505: begin if(four_bit_hash == 0) next_state = 506; else  next_state = 2000;  end 
506: begin if(four_bit_hash == 0) next_state = 507; else  next_state = 2000;  end 
507: begin if(four_bit_hash == 0) next_state = 508; else  next_state = 2000;  end 
508: begin if(four_bit_hash == 0) next_state = 509; else  next_state = 2000;  end 
509: begin if(four_bit_hash == 0) next_state = 510; else  next_state = 2000;  end 
510: begin if(four_bit_hash == 0) next_state = 511; else  next_state = 2000;  end 
511: begin if(four_bit_hash == 0) next_state = 512; else  next_state = 2000;  end 
512: begin if(four_bit_hash == 0) next_state = 513; else  next_state = 2000;  end 
513: begin if(four_bit_hash == 0) next_state = 514; else  next_state = 2000;  end 
514: begin if(four_bit_hash == 0) next_state = 515; else  next_state = 2000;  end 
515: begin if(four_bit_hash == 0) next_state = 516; else  next_state = 2000;  end 
516: begin if(four_bit_hash == 0) next_state = 517; else  next_state = 2000;  end 
517: begin if(four_bit_hash == 0) next_state = 518; else  next_state = 2000;  end 
518: begin if(four_bit_hash == 0) next_state = 519; else  next_state = 2000;  end 
519: begin if(four_bit_hash == 0) next_state = 520; else  next_state = 2000;  end 
520: begin if(four_bit_hash == 0) next_state = 521; else  next_state = 2000;  end 
521: begin if(four_bit_hash == 0) next_state = 522; else  next_state = 2000;  end 
522: begin if(four_bit_hash == 0) next_state = 523; else  next_state = 2000;  end 
523: begin if(four_bit_hash == 0) next_state = 524; else  next_state = 2000;  end 
524: begin if(four_bit_hash == 0) next_state = 525; else  next_state = 2000;  end 
525: begin if(four_bit_hash == 0) next_state = 526; else  next_state = 2000;  end 
526: begin if(four_bit_hash == 0) next_state = 527; else  next_state = 2000;  end 
527: begin if(four_bit_hash == 0) next_state = 528; else  next_state = 2000;  end 
528: begin if(four_bit_hash == 0) next_state = 529; else  next_state = 2000;  end 
529: begin if(four_bit_hash == 0) next_state = 530; else  next_state = 2000;  end 
530: begin if(four_bit_hash == 0) next_state = 531; else  next_state = 2000;  end 
531: begin if(four_bit_hash == 0) next_state = 532; else  next_state = 2000;  end 
532: begin if(four_bit_hash == 0) next_state = 533; else  next_state = 2000;  end 
533: begin if(four_bit_hash == 0) next_state = 534; else  next_state = 2000;  end 
534: begin if(four_bit_hash == 0) next_state = 535; else  next_state = 2000;  end 
535: begin if(four_bit_hash == 0) next_state = 536; else  next_state = 2000;  end 
536: begin if(four_bit_hash == 0) next_state = 537; else  next_state = 2000;  end 
537: begin if(four_bit_hash == 0) next_state = 538; else  next_state = 2000;  end 
538: begin if(four_bit_hash == 0) next_state = 539; else  next_state = 2000;  end 
539: begin if(four_bit_hash == 0) next_state = 540; else  next_state = 2000;  end 
540: begin if(four_bit_hash == 0) next_state = 541; else  next_state = 2000;  end 
541: begin if(four_bit_hash == 0) next_state = 542; else  next_state = 2000;  end 
542: begin if(four_bit_hash == 0) next_state = 543; else  next_state = 2000;  end 
543: begin if(four_bit_hash == 0) next_state = 544; else  next_state = 2000;  end 
544: begin if(four_bit_hash == 0) next_state = 545; else  next_state = 2000;  end 
545: begin if(four_bit_hash == 0) next_state = 546; else  next_state = 2000;  end 
546: begin if(four_bit_hash == 0) next_state = 547; else  next_state = 2000;  end 
547: begin if(four_bit_hash == 0) next_state = 548; else  next_state = 2000;  end 
548: begin if(four_bit_hash == 0) next_state = 549; else  next_state = 2000;  end 
549: begin if(four_bit_hash == 0) next_state = 550; else  next_state = 2000;  end 
550: begin if(four_bit_hash == 0) next_state = 551; else  next_state = 2000;  end 
551: begin if(four_bit_hash == 0) next_state = 552; else  next_state = 2000;  end 
552: begin if(four_bit_hash == 0) next_state = 553; else  next_state = 2000;  end 
553: begin if(four_bit_hash == 0) next_state = 554; else  next_state = 2000;  end 
554: begin if(four_bit_hash == 0) next_state = 555; else  next_state = 2000;  end 
555: begin if(four_bit_hash == 0) next_state = 556; else  next_state = 2000;  end 
556: begin if(four_bit_hash == 0) next_state = 557; else  next_state = 2000;  end 
557: begin if(four_bit_hash == 0) next_state = 558; else  next_state = 2000;  end 
558: begin if(four_bit_hash == 0) next_state = 559; else  next_state = 2000;  end 
559: begin if(four_bit_hash == 0) next_state = 560; else  next_state = 2000;  end 
560: begin if(four_bit_hash == 0) next_state = 561; else  next_state = 2000;  end 
561: begin if(four_bit_hash == 0) next_state = 562; else  next_state = 2000;  end 
562: begin if(four_bit_hash == 0) next_state = 563; else  next_state = 2000;  end 
563: begin if(four_bit_hash == 0) next_state = 564; else  next_state = 2000;  end 
564: begin if(four_bit_hash == 0) next_state = 565; else  next_state = 2000;  end 
565: begin if(four_bit_hash == 0) next_state = 566; else  next_state = 2000;  end 
566: begin if(four_bit_hash == 0) next_state = 567; else  next_state = 2000;  end 
567: begin if(four_bit_hash == 0) next_state = 568; else  next_state = 2000;  end 
568: begin if(four_bit_hash == 0) next_state = 569; else  next_state = 2000;  end 
569: begin if(four_bit_hash == 0) next_state = 570; else  next_state = 2000;  end 
570: begin if(four_bit_hash == 0) next_state = 571; else  next_state = 2000;  end 
571: begin if(four_bit_hash == 0) next_state = 572; else  next_state = 2000;  end 
572: begin if(four_bit_hash == 0) next_state = 573; else  next_state = 2000;  end 
573: begin if(four_bit_hash == 0) next_state = 574; else  next_state = 2000;  end 
574: begin if(four_bit_hash == 0) next_state = 575; else  next_state = 2000;  end 
575: begin if(four_bit_hash == 0) next_state = 576; else  next_state = 2000;  end 
576: begin if(four_bit_hash == 0) next_state = 577; else  next_state = 2000;  end 
577: begin if(four_bit_hash == 0) next_state = 578; else  next_state = 2000;  end 
578: begin if(four_bit_hash == 0) next_state = 579; else  next_state = 2000;  end 
579: begin if(four_bit_hash == 0) next_state = 580; else  next_state = 2000;  end 
580: begin if(four_bit_hash == 0) next_state = 581; else  next_state = 2000;  end 
581: begin if(four_bit_hash == 0) next_state = 582; else  next_state = 2000;  end 
582: begin if(four_bit_hash == 0) next_state = 583; else  next_state = 2000;  end 
583: begin if(four_bit_hash == 0) next_state = 584; else  next_state = 2000;  end 
584: begin if(four_bit_hash == 0) next_state = 585; else  next_state = 2000;  end 
585: begin if(four_bit_hash == 0) next_state = 586; else  next_state = 2000;  end 
586: begin if(four_bit_hash == 0) next_state = 587; else  next_state = 2000;  end 
587: begin if(four_bit_hash == 0) next_state = 588; else  next_state = 2000;  end 
588: begin if(four_bit_hash == 0) next_state = 589; else  next_state = 2000;  end 
589: begin if(four_bit_hash == 0) next_state = 590; else  next_state = 2000;  end 
590: begin if(four_bit_hash == 0) next_state = 591; else  next_state = 2000;  end 
591: begin if(four_bit_hash == 0) next_state = 592; else  next_state = 2000;  end 
592: begin if(four_bit_hash == 0) next_state = 593; else  next_state = 2000;  end 
593: begin if(four_bit_hash == 0) next_state = 594; else  next_state = 2000;  end 
594: begin if(four_bit_hash == 0) next_state = 595; else  next_state = 2000;  end 
595: begin if(four_bit_hash == 0) next_state = 596; else  next_state = 2000;  end 
596: begin if(four_bit_hash == 0) next_state = 597; else  next_state = 2000;  end 
597: begin if(four_bit_hash == 0) next_state = 598; else  next_state = 2000;  end 
598: begin if(four_bit_hash == 0) next_state = 599; else  next_state = 2000;  end 
599: begin if(four_bit_hash == 0) next_state = 600; else  next_state = 2000;  end 
600: begin if(four_bit_hash == 0) next_state = 601; else  next_state = 2000;  end 
601: begin if(four_bit_hash == 0) next_state = 602; else  next_state = 2000;  end 
602: begin if(four_bit_hash == 0) next_state = 603; else  next_state = 2000;  end 
603: begin if(four_bit_hash == 0) next_state = 604; else  next_state = 2000;  end 
604: begin if(four_bit_hash == 0) next_state = 605; else  next_state = 2000;  end 
605: begin if(four_bit_hash == 0) next_state = 606; else  next_state = 2000;  end 
606: begin if(four_bit_hash == 0) next_state = 607; else  next_state = 2000;  end 
607: begin if(four_bit_hash == 0) next_state = 608; else  next_state = 2000;  end 
608: begin if(four_bit_hash == 0) next_state = 609; else  next_state = 2000;  end 
609: begin if(four_bit_hash == 0) next_state = 610; else  next_state = 2000;  end 
610: begin if(four_bit_hash == 0) next_state = 611; else  next_state = 2000;  end 
611: begin if(four_bit_hash == 0) next_state = 612; else  next_state = 2000;  end 
612: begin if(four_bit_hash == 0) next_state = 613; else  next_state = 2000;  end 
613: begin if(four_bit_hash == 0) next_state = 614; else  next_state = 2000;  end 
614: begin if(four_bit_hash == 0) next_state = 615; else  next_state = 2000;  end 
615: begin if(four_bit_hash == 0) next_state = 616; else  next_state = 2000;  end 
616: begin if(four_bit_hash == 0) next_state = 617; else  next_state = 2000;  end 
617: begin if(four_bit_hash == 0) next_state = 618; else  next_state = 2000;  end 
618: begin if(four_bit_hash == 0) next_state = 619; else  next_state = 2000;  end 
619: begin if(four_bit_hash == 0) next_state = 620; else  next_state = 2000;  end 
620: begin if(four_bit_hash == 0) next_state = 621; else  next_state = 2000;  end 
621: begin if(four_bit_hash == 0) next_state = 622; else  next_state = 2000;  end 
622: begin if(four_bit_hash == 0) next_state = 623; else  next_state = 2000;  end 
623: begin if(four_bit_hash == 0) next_state = 624; else  next_state = 2000;  end 
624: begin if(four_bit_hash == 0) next_state = 625; else  next_state = 2000;  end 
625: begin if(four_bit_hash == 0) next_state = 626; else  next_state = 2000;  end 
626: begin if(four_bit_hash == 0) next_state = 627; else  next_state = 2000;  end 
627: begin if(four_bit_hash == 0) next_state = 628; else  next_state = 2000;  end 
628: begin if(four_bit_hash == 0) next_state = 629; else  next_state = 2000;  end 
629: begin if(four_bit_hash == 0) next_state = 630; else  next_state = 2000;  end 
630: begin if(four_bit_hash == 0) next_state = 631; else  next_state = 2000;  end 
631: begin if(four_bit_hash == 0) next_state = 632; else  next_state = 2000;  end 
632: begin if(four_bit_hash == 0) next_state = 633; else  next_state = 2000;  end 
633: begin if(four_bit_hash == 0) next_state = 634; else  next_state = 2000;  end 
634: begin if(four_bit_hash == 0) next_state = 635; else  next_state = 2000;  end 
635: begin if(four_bit_hash == 0) next_state = 636; else  next_state = 2000;  end 
636: begin if(four_bit_hash == 0) next_state = 637; else  next_state = 2000;  end 
637: begin if(four_bit_hash == 0) next_state = 638; else  next_state = 2000;  end 
638: begin if(four_bit_hash == 0) next_state = 639; else  next_state = 2000;  end 
639: begin if(four_bit_hash == 0) next_state = 640; else  next_state = 2000;  end 
640: begin if(four_bit_hash == 0) next_state = 641; else  next_state = 2000;  end 
641: begin if(four_bit_hash == 0) next_state = 642; else  next_state = 2000;  end 
642: begin if(four_bit_hash == 0) next_state = 643; else  next_state = 2000;  end 
643: begin if(four_bit_hash == 0) next_state = 644; else  next_state = 2000;  end 
644: begin if(four_bit_hash == 0) next_state = 645; else  next_state = 2000;  end 
645: begin if(four_bit_hash == 0) next_state = 646; else  next_state = 2000;  end 
646: begin if(four_bit_hash == 0) next_state = 647; else  next_state = 2000;  end 
647: begin if(four_bit_hash == 0) next_state = 648; else  next_state = 2000;  end 
648: begin if(four_bit_hash == 0) next_state = 649; else  next_state = 2000;  end 
649: begin if(four_bit_hash == 0) next_state = 650; else  next_state = 2000;  end 
650: begin if(four_bit_hash == 0) next_state = 651; else  next_state = 2000;  end 
651: begin if(four_bit_hash == 0) next_state = 652; else  next_state = 2000;  end 
652: begin if(four_bit_hash == 0) next_state = 653; else  next_state = 2000;  end 
653: begin if(four_bit_hash == 0) next_state = 654; else  next_state = 2000;  end 
654: begin if(four_bit_hash == 0) next_state = 655; else  next_state = 2000;  end 
655: begin if(four_bit_hash == 0) next_state = 656; else  next_state = 2000;  end 
656: begin if(four_bit_hash == 0) next_state = 657; else  next_state = 2000;  end 
657: begin if(four_bit_hash == 0) next_state = 658; else  next_state = 2000;  end 
658: begin if(four_bit_hash == 0) next_state = 659; else  next_state = 2000;  end 
659: begin if(four_bit_hash == 0) next_state = 660; else  next_state = 2000;  end 
660: begin if(four_bit_hash == 0) next_state = 661; else  next_state = 2000;  end 
661: begin if(four_bit_hash == 0) next_state = 662; else  next_state = 2000;  end 
662: begin if(four_bit_hash == 0) next_state = 663; else  next_state = 2000;  end 
663: begin if(four_bit_hash == 0) next_state = 664; else  next_state = 2000;  end 
664: begin if(four_bit_hash == 0) next_state = 665; else  next_state = 2000;  end 
665: begin if(four_bit_hash == 0) next_state = 666; else  next_state = 2000;  end 
666: begin if(four_bit_hash == 0) next_state = 667; else  next_state = 2000;  end 
667: begin if(four_bit_hash == 0) next_state = 668; else  next_state = 2000;  end 
668: begin if(four_bit_hash == 0) next_state = 669; else  next_state = 2000;  end 
669: begin if(four_bit_hash == 0) next_state = 670; else  next_state = 2000;  end 
670: begin if(four_bit_hash == 0) next_state = 671; else  next_state = 2000;  end 
671: begin if(four_bit_hash == 0) next_state = 672; else  next_state = 2000;  end 
672: begin if(four_bit_hash == 0) next_state = 673; else  next_state = 2000;  end 
673: begin if(four_bit_hash == 0) next_state = 674; else  next_state = 2000;  end 
674: begin if(four_bit_hash == 0) next_state = 675; else  next_state = 2000;  end 
675: begin if(four_bit_hash == 0) next_state = 676; else  next_state = 2000;  end 
676: begin if(four_bit_hash == 0) next_state = 677; else  next_state = 2000;  end 
677: begin if(four_bit_hash == 0) next_state = 678; else  next_state = 2000;  end 
678: begin if(four_bit_hash == 0) next_state = 679; else  next_state = 2000;  end 
679: begin if(four_bit_hash == 0) next_state = 680; else  next_state = 2000;  end 
680: begin if(four_bit_hash == 0) next_state = 681; else  next_state = 2000;  end 
681: begin if(four_bit_hash == 0) next_state = 682; else  next_state = 2000;  end 
682: begin if(four_bit_hash == 0) next_state = 683; else  next_state = 2000;  end 
683: begin if(four_bit_hash == 0) next_state = 684; else  next_state = 2000;  end 
684: begin if(four_bit_hash == 0) next_state = 685; else  next_state = 2000;  end 
685: begin if(four_bit_hash == 0) next_state = 686; else  next_state = 2000;  end 
686: begin if(four_bit_hash == 0) next_state = 687; else  next_state = 2000;  end 
687: begin if(four_bit_hash == 0) next_state = 688; else  next_state = 2000;  end 
688: begin if(four_bit_hash == 0) next_state = 689; else  next_state = 2000;  end 
689: begin if(four_bit_hash == 0) next_state = 690; else  next_state = 2000;  end 
690: begin if(four_bit_hash == 0) next_state = 691; else  next_state = 2000;  end 
691: begin if(four_bit_hash == 0) next_state = 692; else  next_state = 2000;  end 
692: begin if(four_bit_hash == 0) next_state = 693; else  next_state = 2000;  end 
693: begin if(four_bit_hash == 0) next_state = 694; else  next_state = 2000;  end 
694: begin if(four_bit_hash == 0) next_state = 695; else  next_state = 2000;  end 
695: begin if(four_bit_hash == 0) next_state = 696; else  next_state = 2000;  end 
696: begin if(four_bit_hash == 0) next_state = 697; else  next_state = 2000;  end 
697: begin if(four_bit_hash == 0) next_state = 698; else  next_state = 2000;  end 
698: begin if(four_bit_hash == 0) next_state = 699; else  next_state = 2000;  end 
699: begin if(four_bit_hash == 0) next_state = 700; else  next_state = 2000;  end 
700: begin if(four_bit_hash == 0) next_state = 701; else  next_state = 2000;  end 
701: begin if(four_bit_hash == 0) next_state = 702; else  next_state = 2000;  end 
702: begin if(four_bit_hash == 0) next_state = 703; else  next_state = 2000;  end 
703: begin if(four_bit_hash == 0) next_state = 704; else  next_state = 2000;  end 
704: begin if(four_bit_hash == 0) next_state = 705; else  next_state = 2000;  end 
705: begin if(four_bit_hash == 0) next_state = 706; else  next_state = 2000;  end 
706: begin if(four_bit_hash == 0) next_state = 707; else  next_state = 2000;  end 
707: begin if(four_bit_hash == 0) next_state = 708; else  next_state = 2000;  end 
708: begin if(four_bit_hash == 0) next_state = 709; else  next_state = 2000;  end 
709: begin if(four_bit_hash == 0) next_state = 710; else  next_state = 2000;  end 
710: begin if(four_bit_hash == 0) next_state = 711; else  next_state = 2000;  end 
711: begin if(four_bit_hash == 0) next_state = 712; else  next_state = 2000;  end 
712: begin if(four_bit_hash == 0) next_state = 713; else  next_state = 2000;  end 
713: begin if(four_bit_hash == 0) next_state = 714; else  next_state = 2000;  end 
714: begin if(four_bit_hash == 0) next_state = 715; else  next_state = 2000;  end 
715: begin if(four_bit_hash == 0) next_state = 716; else  next_state = 2000;  end 
716: begin if(four_bit_hash == 0) next_state = 717; else  next_state = 2000;  end 
717: begin if(four_bit_hash == 0) next_state = 718; else  next_state = 2000;  end 
718: begin if(four_bit_hash == 0) next_state = 719; else  next_state = 2000;  end 
719: begin if(four_bit_hash == 0) next_state = 720; else  next_state = 2000;  end 
720: begin if(four_bit_hash == 0) next_state = 721; else  next_state = 2000;  end 
721: begin if(four_bit_hash == 0) next_state = 722; else  next_state = 2000;  end 
722: begin if(four_bit_hash == 0) next_state = 723; else  next_state = 2000;  end 
723: begin if(four_bit_hash == 0) next_state = 724; else  next_state = 2000;  end 
724: begin if(four_bit_hash == 0) next_state = 725; else  next_state = 2000;  end 
725: begin if(four_bit_hash == 0) next_state = 726; else  next_state = 2000;  end 
726: begin if(four_bit_hash == 0) next_state = 727; else  next_state = 2000;  end 
727: begin if(four_bit_hash == 0) next_state = 728; else  next_state = 2000;  end 
728: begin if(four_bit_hash == 0) next_state = 729; else  next_state = 2000;  end 
729: begin if(four_bit_hash == 0) next_state = 730; else  next_state = 2000;  end 
730: begin if(four_bit_hash == 0) next_state = 731; else  next_state = 2000;  end 
731: begin if(four_bit_hash == 0) next_state = 732; else  next_state = 2000;  end 
732: begin if(four_bit_hash == 0) next_state = 733; else  next_state = 2000;  end 
733: begin if(four_bit_hash == 0) next_state = 734; else  next_state = 2000;  end 
734: begin if(four_bit_hash == 0) next_state = 735; else  next_state = 2000;  end 
735: begin if(four_bit_hash == 0) next_state = 736; else  next_state = 2000;  end 
736: begin if(four_bit_hash == 0) next_state = 737; else  next_state = 2000;  end 
737: begin if(four_bit_hash == 0) next_state = 738; else  next_state = 2000;  end 
738: begin if(four_bit_hash == 0) next_state = 739; else  next_state = 2000;  end 
739: begin if(four_bit_hash == 0) next_state = 740; else  next_state = 2000;  end 
740: begin if(four_bit_hash == 0) next_state = 741; else  next_state = 2000;  end 
741: begin if(four_bit_hash == 0) next_state = 742; else  next_state = 2000;  end 
742: begin if(four_bit_hash == 0) next_state = 743; else  next_state = 2000;  end 
743: begin if(four_bit_hash == 0) next_state = 744; else  next_state = 2000;  end 
744: begin if(four_bit_hash == 0) next_state = 745; else  next_state = 2000;  end 
745: begin if(four_bit_hash == 0) next_state = 746; else  next_state = 2000;  end 
746: begin if(four_bit_hash == 0) next_state = 747; else  next_state = 2000;  end 
747: begin if(four_bit_hash == 0) next_state = 748; else  next_state = 2000;  end 
748: begin if(four_bit_hash == 0) next_state = 749; else  next_state = 2000;  end 
749: begin if(four_bit_hash == 0) next_state = 750; else  next_state = 2000;  end 
750: begin if(four_bit_hash == 0) next_state = 751; else  next_state = 2000;  end 
751: begin if(four_bit_hash == 0) next_state = 752; else  next_state = 2000;  end 
752: begin if(four_bit_hash == 0) next_state = 753; else  next_state = 2000;  end 
753: begin if(four_bit_hash == 0) next_state = 754; else  next_state = 2000;  end 
754: begin if(four_bit_hash == 0) next_state = 755; else  next_state = 2000;  end 
755: begin if(four_bit_hash == 0) next_state = 756; else  next_state = 2000;  end 
756: begin if(four_bit_hash == 0) next_state = 757; else  next_state = 2000;  end 
757: begin if(four_bit_hash == 0) next_state = 758; else  next_state = 2000;  end 
758: begin if(four_bit_hash == 0) next_state = 759; else  next_state = 2000;  end 
759: begin if(four_bit_hash == 0) next_state = 760; else  next_state = 2000;  end 
760: begin if(four_bit_hash == 0) next_state = 761; else  next_state = 2000;  end 
761: begin if(four_bit_hash == 0) next_state = 762; else  next_state = 2000;  end 
762: begin if(four_bit_hash == 0) next_state = 763; else  next_state = 2000;  end 
763: begin if(four_bit_hash == 0) next_state = 764; else  next_state = 2000;  end 
764: begin if(four_bit_hash == 0) next_state = 765; else  next_state = 2000;  end 
765: begin if(four_bit_hash == 0) next_state = 766; else  next_state = 2000;  end 
766: begin if(four_bit_hash == 0) next_state = 767; else  next_state = 2000;  end 
767: begin if(four_bit_hash == 0) next_state = 768; else  next_state = 2000;  end 
768: begin if(four_bit_hash == 0) next_state = 769; else  next_state = 2000;  end 
769: begin if(four_bit_hash == 0) next_state = 770; else  next_state = 2000;  end 
770: begin if(four_bit_hash == 0) next_state = 771; else  next_state = 2000;  end 
771: begin if(four_bit_hash == 0) next_state = 772; else  next_state = 2000;  end 
772: begin if(four_bit_hash == 0) next_state = 773; else  next_state = 2000;  end 
773: begin if(four_bit_hash == 0) next_state = 774; else  next_state = 2000;  end 
774: begin if(four_bit_hash == 0) next_state = 775; else  next_state = 2000;  end 
775: begin if(four_bit_hash == 0) next_state = 776; else  next_state = 2000;  end 
776: begin if(four_bit_hash == 0) next_state = 777; else  next_state = 2000;  end 
777: begin if(four_bit_hash == 0) next_state = 778; else  next_state = 2000;  end 
778: begin if(four_bit_hash == 0) next_state = 779; else  next_state = 2000;  end 
779: begin if(four_bit_hash == 0) next_state = 780; else  next_state = 2000;  end 
780: begin if(four_bit_hash == 0) next_state = 781; else  next_state = 2000;  end 
781: begin if(four_bit_hash == 0) next_state = 782; else  next_state = 2000;  end 
782: begin if(four_bit_hash == 0) next_state = 783; else  next_state = 2000;  end 
783: begin if(four_bit_hash == 0) next_state = 784; else  next_state = 2000;  end 
784: begin if(four_bit_hash == 0) next_state = 785; else  next_state = 2000;  end 
785: begin if(four_bit_hash == 0) next_state = 786; else  next_state = 2000;  end 
786: begin if(four_bit_hash == 0) next_state = 787; else  next_state = 2000;  end 
787: begin if(four_bit_hash == 0) next_state = 788; else  next_state = 2000;  end 
788: begin if(four_bit_hash == 0) next_state = 789; else  next_state = 2000;  end 
789: begin if(four_bit_hash == 0) next_state = 790; else  next_state = 2000;  end 
790: begin if(four_bit_hash == 0) next_state = 791; else  next_state = 2000;  end 
791: begin if(four_bit_hash == 0) next_state = 792; else  next_state = 2000;  end 
792: begin if(four_bit_hash == 0) next_state = 793; else  next_state = 2000;  end 
793: begin if(four_bit_hash == 0) next_state = 794; else  next_state = 2000;  end 
794: begin if(four_bit_hash == 0) next_state = 795; else  next_state = 2000;  end 
795: begin if(four_bit_hash == 0) next_state = 796; else  next_state = 2000;  end 
796: begin if(four_bit_hash == 0) next_state = 797; else  next_state = 2000;  end 
797: begin if(four_bit_hash == 0) next_state = 798; else  next_state = 2000;  end 
798: begin if(four_bit_hash == 0) next_state = 799; else  next_state = 2000;  end 
799: begin if(four_bit_hash == 0) next_state = 800; else  next_state = 2000;  end 
800: begin if(four_bit_hash == 0) next_state = 801; else  next_state = 2000;  end 
801: begin if(four_bit_hash == 0) next_state = 802; else  next_state = 2000;  end 
802: begin if(four_bit_hash == 0) next_state = 803; else  next_state = 2000;  end 
803: begin if(four_bit_hash == 0) next_state = 804; else  next_state = 2000;  end 
804: begin if(four_bit_hash == 0) next_state = 805; else  next_state = 2000;  end 
805: begin if(four_bit_hash == 0) next_state = 806; else  next_state = 2000;  end 
806: begin if(four_bit_hash == 0) next_state = 807; else  next_state = 2000;  end 
807: begin if(four_bit_hash == 0) next_state = 808; else  next_state = 2000;  end 
808: begin if(four_bit_hash == 0) next_state = 809; else  next_state = 2000;  end 
809: begin if(four_bit_hash == 0) next_state = 810; else  next_state = 2000;  end 
810: begin if(four_bit_hash == 0) next_state = 811; else  next_state = 2000;  end 
811: begin if(four_bit_hash == 0) next_state = 812; else  next_state = 2000;  end 
812: begin if(four_bit_hash == 0) next_state = 813; else  next_state = 2000;  end 
813: begin if(four_bit_hash == 0) next_state = 814; else  next_state = 2000;  end 
814: begin if(four_bit_hash == 0) next_state = 815; else  next_state = 2000;  end 
815: begin if(four_bit_hash == 0) next_state = 816; else  next_state = 2000;  end 
816: begin if(four_bit_hash == 0) next_state = 817; else  next_state = 2000;  end 
817: begin if(four_bit_hash == 0) next_state = 818; else  next_state = 2000;  end 
818: begin if(four_bit_hash == 0) next_state = 819; else  next_state = 2000;  end 
819: begin if(four_bit_hash == 0) next_state = 820; else  next_state = 2000;  end 
820: begin if(four_bit_hash == 0) next_state = 821; else  next_state = 2000;  end 
821: begin if(four_bit_hash == 0) next_state = 822; else  next_state = 2000;  end 
822: begin if(four_bit_hash == 0) next_state = 823; else  next_state = 2000;  end 
823: begin if(four_bit_hash == 0) next_state = 824; else  next_state = 2000;  end 
824: begin if(four_bit_hash == 0) next_state = 825; else  next_state = 2000;  end 
825: begin if(four_bit_hash == 0) next_state = 826; else  next_state = 2000;  end 
826: begin if(four_bit_hash == 0) next_state = 827; else  next_state = 2000;  end 
827: begin if(four_bit_hash == 0) next_state = 828; else  next_state = 2000;  end 
828: begin if(four_bit_hash == 0) next_state = 829; else  next_state = 2000;  end 
829: begin if(four_bit_hash == 0) next_state = 830; else  next_state = 2000;  end 
830: begin if(four_bit_hash == 0) next_state = 831; else  next_state = 2000;  end 
831: begin if(four_bit_hash == 0) next_state = 832; else  next_state = 2000;  end 
832: begin if(four_bit_hash == 0) next_state = 833; else  next_state = 2000;  end 
833: begin if(four_bit_hash == 0) next_state = 834; else  next_state = 2000;  end 
834: begin if(four_bit_hash == 0) next_state = 835; else  next_state = 2000;  end 
835: begin if(four_bit_hash == 0) next_state = 836; else  next_state = 2000;  end 
836: begin if(four_bit_hash == 0) next_state = 837; else  next_state = 2000;  end 
837: begin if(four_bit_hash == 0) next_state = 838; else  next_state = 2000;  end 
838: begin if(four_bit_hash == 0) next_state = 839; else  next_state = 2000;  end 
839: begin if(four_bit_hash == 0) next_state = 840; else  next_state = 2000;  end 
840: begin if(four_bit_hash == 0) next_state = 841; else  next_state = 2000;  end 
841: begin if(four_bit_hash == 0) next_state = 842; else  next_state = 2000;  end 
842: begin if(four_bit_hash == 0) next_state = 843; else  next_state = 2000;  end 
843: begin if(four_bit_hash == 0) next_state = 844; else  next_state = 2000;  end 
844: begin if(four_bit_hash == 0) next_state = 845; else  next_state = 2000;  end 
845: begin if(four_bit_hash == 0) next_state = 846; else  next_state = 2000;  end 
846: begin if(four_bit_hash == 0) next_state = 847; else  next_state = 2000;  end 
847: begin if(four_bit_hash == 0) next_state = 848; else  next_state = 2000;  end 
848: begin if(four_bit_hash == 0) next_state = 849; else  next_state = 2000;  end 
849: begin if(four_bit_hash == 0) next_state = 850; else  next_state = 2000;  end 
850: begin if(four_bit_hash == 0) next_state = 851; else  next_state = 2000;  end 
851: begin if(four_bit_hash == 0) next_state = 852; else  next_state = 2000;  end 
852: begin if(four_bit_hash == 0) next_state = 853; else  next_state = 2000;  end 
853: begin if(four_bit_hash == 0) next_state = 854; else  next_state = 2000;  end 
854: begin if(four_bit_hash == 0) next_state = 855; else  next_state = 2000;  end 
855: begin if(four_bit_hash == 0) next_state = 856; else  next_state = 2000;  end 
856: begin if(four_bit_hash == 0) next_state = 857; else  next_state = 2000;  end 
857: begin if(four_bit_hash == 0) next_state = 858; else  next_state = 2000;  end 
858: begin if(four_bit_hash == 0) next_state = 859; else  next_state = 2000;  end 
859: begin if(four_bit_hash == 0) next_state = 860; else  next_state = 2000;  end 
860: begin if(four_bit_hash == 0) next_state = 861; else  next_state = 2000;  end 
861: begin if(four_bit_hash == 0) next_state = 862; else  next_state = 2000;  end 
862: begin if(four_bit_hash == 0) next_state = 863; else  next_state = 2000;  end 
863: begin if(four_bit_hash == 0) next_state = 864; else  next_state = 2000;  end 
864: begin if(four_bit_hash == 0) next_state = 865; else  next_state = 2000;  end 
865: begin if(four_bit_hash == 0) next_state = 866; else  next_state = 2000;  end 
866: begin if(four_bit_hash == 0) next_state = 867; else  next_state = 2000;  end 
867: begin if(four_bit_hash == 0) next_state = 868; else  next_state = 2000;  end 
868: begin if(four_bit_hash == 0) next_state = 869; else  next_state = 2000;  end 
869: begin if(four_bit_hash == 0) next_state = 870; else  next_state = 2000;  end 
870: begin if(four_bit_hash == 0) next_state = 871; else  next_state = 2000;  end 
871: begin if(four_bit_hash == 0) next_state = 872; else  next_state = 2000;  end 
872: begin if(four_bit_hash == 0) next_state = 873; else  next_state = 2000;  end 
873: begin if(four_bit_hash == 0) next_state = 874; else  next_state = 2000;  end 
874: begin if(four_bit_hash == 0) next_state = 875; else  next_state = 2000;  end 
875: begin if(four_bit_hash == 0) next_state = 876; else  next_state = 2000;  end 
876: begin if(four_bit_hash == 0) next_state = 877; else  next_state = 2000;  end 
877: begin if(four_bit_hash == 0) next_state = 878; else  next_state = 2000;  end 
878: begin if(four_bit_hash == 0) next_state = 879; else  next_state = 2000;  end 
879: begin if(four_bit_hash == 0) next_state = 880; else  next_state = 2000;  end 
880: begin if(four_bit_hash == 0) next_state = 881; else  next_state = 2000;  end 
881: begin if(four_bit_hash == 0) next_state = 882; else  next_state = 2000;  end 
882: begin if(four_bit_hash == 0) next_state = 883; else  next_state = 2000;  end 
883: begin if(four_bit_hash == 0) next_state = 884; else  next_state = 2000;  end 
884: begin if(four_bit_hash == 0) next_state = 885; else  next_state = 2000;  end 
885: begin if(four_bit_hash == 0) next_state = 886; else  next_state = 2000;  end 
886: begin if(four_bit_hash == 0) next_state = 887; else  next_state = 2000;  end 
887: begin if(four_bit_hash == 0) next_state = 888; else  next_state = 2000;  end 
888: begin if(four_bit_hash == 0) next_state = 889; else  next_state = 2000;  end 
889: begin if(four_bit_hash == 0) next_state = 890; else  next_state = 2000;  end 
890: begin if(four_bit_hash == 0) next_state = 891; else  next_state = 2000;  end 
891: begin if(four_bit_hash == 0) next_state = 892; else  next_state = 2000;  end 
892: begin if(four_bit_hash == 0) next_state = 893; else  next_state = 2000;  end 
893: begin if(four_bit_hash == 0) next_state = 894; else  next_state = 2000;  end 
894: begin if(four_bit_hash == 0) next_state = 895; else  next_state = 2000;  end 
895: begin if(four_bit_hash == 0) next_state = 896; else  next_state = 2000;  end 
896: begin if(four_bit_hash == 0) next_state = 897; else  next_state = 2000;  end 
897: begin if(four_bit_hash == 0) next_state = 898; else  next_state = 2000;  end 
898: begin if(four_bit_hash == 0) next_state = 899; else  next_state = 2000;  end 
899: begin if(four_bit_hash == 0) next_state = 900; else  next_state = 2000;  end 
900: begin if(four_bit_hash == 0) next_state = 901; else  next_state = 2000;  end 
901: begin if(four_bit_hash == 0) next_state = 902; else  next_state = 2000;  end 
902: begin if(four_bit_hash == 0) next_state = 903; else  next_state = 2000;  end 
903: begin if(four_bit_hash == 0) next_state = 904; else  next_state = 2000;  end 
904: begin if(four_bit_hash == 0) next_state = 905; else  next_state = 2000;  end 
905: begin if(four_bit_hash == 0) next_state = 906; else  next_state = 2000;  end 
906: begin if(four_bit_hash == 0) next_state = 907; else  next_state = 2000;  end 
907: begin if(four_bit_hash == 0) next_state = 908; else  next_state = 2000;  end 
908: begin if(four_bit_hash == 0) next_state = 909; else  next_state = 2000;  end 
909: begin if(four_bit_hash == 0) next_state = 910; else  next_state = 2000;  end 
910: begin if(four_bit_hash == 0) next_state = 911; else  next_state = 2000;  end 
911: begin if(four_bit_hash == 0) next_state = 912; else  next_state = 2000;  end 
912: begin if(four_bit_hash == 0) next_state = 913; else  next_state = 2000;  end 
913: begin if(four_bit_hash == 0) next_state = 914; else  next_state = 2000;  end 
914: begin if(four_bit_hash == 0) next_state = 915; else  next_state = 2000;  end 
915: begin if(four_bit_hash == 0) next_state = 916; else  next_state = 2000;  end 
916: begin if(four_bit_hash == 0) next_state = 917; else  next_state = 2000;  end 
917: begin if(four_bit_hash == 0) next_state = 918; else  next_state = 2000;  end 
918: begin if(four_bit_hash == 0) next_state = 919; else  next_state = 2000;  end 
919: begin if(four_bit_hash == 0) next_state = 920; else  next_state = 2000;  end 
920: begin if(four_bit_hash == 0) next_state = 921; else  next_state = 2000;  end 
921: begin if(four_bit_hash == 0) next_state = 922; else  next_state = 2000;  end 
922: begin if(four_bit_hash == 0) next_state = 923; else  next_state = 2000;  end 
923: begin if(four_bit_hash == 0) next_state = 924; else  next_state = 2000;  end 
924: begin if(four_bit_hash == 0) next_state = 925; else  next_state = 2000;  end 
925: begin if(four_bit_hash == 0) next_state = 926; else  next_state = 2000;  end 
926: begin if(four_bit_hash == 0) next_state = 927; else  next_state = 2000;  end 
927: begin if(four_bit_hash == 0) next_state = 928; else  next_state = 2000;  end 
928: begin if(four_bit_hash == 0) next_state = 929; else  next_state = 2000;  end 
929: begin if(four_bit_hash == 0) next_state = 930; else  next_state = 2000;  end 
930: begin if(four_bit_hash == 0) next_state = 931; else  next_state = 2000;  end 
931: begin if(four_bit_hash == 0) next_state = 932; else  next_state = 2000;  end 
932: begin if(four_bit_hash == 0) next_state = 933; else  next_state = 2000;  end 
933: begin if(four_bit_hash == 0) next_state = 934; else  next_state = 2000;  end 
934: begin if(four_bit_hash == 0) next_state = 935; else  next_state = 2000;  end 
935: begin if(four_bit_hash == 0) next_state = 936; else  next_state = 2000;  end 
936: begin if(four_bit_hash == 0) next_state = 937; else  next_state = 2000;  end 
937: begin if(four_bit_hash == 0) next_state = 938; else  next_state = 2000;  end 
938: begin if(four_bit_hash == 0) next_state = 939; else  next_state = 2000;  end 
939: begin if(four_bit_hash == 0) next_state = 940; else  next_state = 2000;  end 
940: begin if(four_bit_hash == 0) next_state = 941; else  next_state = 2000;  end 
941: begin if(four_bit_hash == 0) next_state = 942; else  next_state = 2000;  end 
942: begin if(four_bit_hash == 0) next_state = 943; else  next_state = 2000;  end 
943: begin if(four_bit_hash == 0) next_state = 944; else  next_state = 2000;  end 
944: begin if(four_bit_hash == 0) next_state = 945; else  next_state = 2000;  end 
945: begin if(four_bit_hash == 0) next_state = 946; else  next_state = 2000;  end 
946: begin if(four_bit_hash == 0) next_state = 947; else  next_state = 2000;  end 
947: begin if(four_bit_hash == 0) next_state = 948; else  next_state = 2000;  end 
948: begin if(four_bit_hash == 0) next_state = 949; else  next_state = 2000;  end 
949: begin if(four_bit_hash == 0) next_state = 950; else  next_state = 2000;  end 
950: begin if(four_bit_hash == 0) next_state = 951; else  next_state = 2000;  end 
951: begin if(four_bit_hash == 0) next_state = 952; else  next_state = 2000;  end 
952: begin if(four_bit_hash == 0) next_state = 953; else  next_state = 2000;  end 
953: begin if(four_bit_hash == 0) next_state = 954; else  next_state = 2000;  end 
954: begin if(four_bit_hash == 0) next_state = 955; else  next_state = 2000;  end 
955: begin if(four_bit_hash == 0) next_state = 956; else  next_state = 2000;  end 
956: begin if(four_bit_hash == 0) next_state = 957; else  next_state = 2000;  end 
957: begin if(four_bit_hash == 0) next_state = 958; else  next_state = 2000;  end 
958: begin if(four_bit_hash == 0) next_state = 959; else  next_state = 2000;  end 
959: begin if(four_bit_hash == 0) next_state = 960; else  next_state = 2000;  end 
960: begin if(four_bit_hash == 0) next_state = 961; else  next_state = 2000;  end 
961: begin if(four_bit_hash == 0) next_state = 962; else  next_state = 2000;  end 
962: begin if(four_bit_hash == 0) next_state = 963; else  next_state = 2000;  end 
963: begin if(four_bit_hash == 0) next_state = 964; else  next_state = 2000;  end 
964: begin if(four_bit_hash == 0) next_state = 965; else  next_state = 2000;  end 
965: begin if(four_bit_hash == 0) next_state = 966; else  next_state = 2000;  end 
966: begin if(four_bit_hash == 0) next_state = 967; else  next_state = 2000;  end 
967: begin if(four_bit_hash == 0) next_state = 968; else  next_state = 2000;  end 
968: begin if(four_bit_hash == 0) next_state = 969; else  next_state = 2000;  end 
969: begin if(four_bit_hash == 0) next_state = 970; else  next_state = 2000;  end 
970: begin if(four_bit_hash == 0) next_state = 971; else  next_state = 2000;  end 
971: begin if(four_bit_hash == 0) next_state = 972; else  next_state = 2000;  end 
972: begin if(four_bit_hash == 0) next_state = 973; else  next_state = 2000;  end 
973: begin if(four_bit_hash == 0) next_state = 974; else  next_state = 2000;  end 
974: begin if(four_bit_hash == 0) next_state = 975; else  next_state = 2000;  end 
975: begin if(four_bit_hash == 0) next_state = 976; else  next_state = 2000;  end 
976: begin if(four_bit_hash == 0) next_state = 977; else  next_state = 2000;  end 
977: begin if(four_bit_hash == 0) next_state = 978; else  next_state = 2000;  end 
978: begin if(four_bit_hash == 0) next_state = 979; else  next_state = 2000;  end 
979: begin if(four_bit_hash == 0) next_state = 980; else  next_state = 2000;  end 
980: begin if(four_bit_hash == 0) next_state = 981; else  next_state = 2000;  end 
981: begin if(four_bit_hash == 0) next_state = 982; else  next_state = 2000;  end 
982: begin if(four_bit_hash == 0) next_state = 983; else  next_state = 2000;  end 
983: begin if(four_bit_hash == 0) next_state = 984; else  next_state = 2000;  end 
984: begin if(four_bit_hash == 0) next_state = 985; else  next_state = 2000;  end 
985: begin if(four_bit_hash == 0) next_state = 986; else  next_state = 2000;  end 
986: begin if(four_bit_hash == 0) next_state = 987; else  next_state = 2000;  end 
987: begin if(four_bit_hash == 0) next_state = 988; else  next_state = 2000;  end 
988: begin if(four_bit_hash == 0) next_state = 989; else  next_state = 2000;  end 
989: begin if(four_bit_hash == 0) next_state = 990; else  next_state = 2000;  end 
990: begin if(four_bit_hash == 0) next_state = 991; else  next_state = 2000;  end 
991: begin if(four_bit_hash == 0) next_state = 992; else  next_state = 2000;  end 
992: begin if(four_bit_hash == 0) next_state = 993; else  next_state = 2000;  end 
993: begin if(four_bit_hash == 0) next_state = 994; else  next_state = 2000;  end 
994: begin if(four_bit_hash == 0) next_state = 995; else  next_state = 2000;  end 
995: begin if(four_bit_hash == 0) next_state = 996; else  next_state = 2000;  end 
996: begin if(four_bit_hash == 0) next_state = 997; else  next_state = 2000;  end 
997: begin if(four_bit_hash == 0) next_state = 998; else  next_state = 2000;  end 
998: begin if(four_bit_hash == 0) next_state = 999; else  next_state = 2000;  end 
999: begin if(four_bit_hash == 0) next_state = 1000; else  next_state = 2000;  end 
1000: begin if(four_bit_hash == 0) next_state = 1001; else  next_state = 2000;  end 
1001: begin if(four_bit_hash == 0) next_state = 1002; else  next_state = 2000;  end 
1002: begin if(four_bit_hash == 0) next_state = 1003; else  next_state = 2000;  end 
1003: begin if(four_bit_hash == 0) next_state = 1004; else  next_state = 2000;  end 
1004: begin if(four_bit_hash == 0) next_state = 1005; else  next_state = 2000;  end 
1005: begin if(four_bit_hash == 0) next_state = 1006; else  next_state = 2000;  end 
1006: begin if(four_bit_hash == 0) next_state = 1007; else  next_state = 2000;  end 
1007: begin if(four_bit_hash == 0) next_state = 1008; else  next_state = 2000;  end 
1008: begin if(four_bit_hash == 0) next_state = 1009; else  next_state = 2000;  end 
1009: begin if(four_bit_hash == 0) next_state = 1010; else  next_state = 2000;  end 
1010: begin if(four_bit_hash == 0) next_state = 1011; else  next_state = 2000;  end 
1011: begin if(four_bit_hash == 0) next_state = 1012; else  next_state = 2000;  end 
1012: begin if(four_bit_hash == 0) next_state = 1013; else  next_state = 2000;  end 
1013: begin if(four_bit_hash == 0) next_state = 1014; else  next_state = 2000;  end 
1014: begin if(four_bit_hash == 0) next_state = 1015; else  next_state = 2000;  end 
1015: begin if(four_bit_hash == 0) next_state = 1016; else  next_state = 2000;  end 
1016: begin if(four_bit_hash == 0) next_state = 1017; else  next_state = 2000;  end 
1017: begin if(four_bit_hash == 0) next_state = 1018; else  next_state = 2000;  end 
1018: begin if(four_bit_hash == 0) next_state = 1019; else  next_state = 2000;  end 
1019: begin if(four_bit_hash == 0) next_state = 1020; else  next_state = 2000;  end 
1020: begin if(four_bit_hash == 0) next_state = 1021; else  next_state = 2000;  end 
1021: begin if(four_bit_hash == 0) next_state = 1022; else  next_state = 2000;  end 
1022: begin if(four_bit_hash == 0) next_state = 1023; else  next_state = 2000;  end 
1023: begin if(four_bit_hash == 0) next_state = 1024; else  next_state = 2000;  end 
1024: begin if(four_bit_hash == 0) next_state = 1025; else  next_state = 2000;  end 
1025: begin if(four_bit_hash == 0) next_state = 1026; else  next_state = 2000;  end 
1026: begin if(four_bit_hash == 0) next_state = 1027; else  next_state = 2000;  end 
1027: begin if(four_bit_hash == 0) next_state = 1028; else  next_state = 2000;  end 
1028: begin if(four_bit_hash == 0) next_state = 1029; else  next_state = 2000;  end 
1029: begin if(four_bit_hash == 0) next_state = 1030; else  next_state = 2000;  end 
1030: begin if(four_bit_hash == 0) next_state = 1031; else  next_state = 2000;  end 
1031: begin if(four_bit_hash == 0) next_state = 1032; else  next_state = 2000;  end 
1032: begin if(four_bit_hash == 0) next_state = 1033; else  next_state = 2000;  end 
1033: begin if(four_bit_hash == 0) next_state = 1034; else  next_state = 2000;  end 
1034: begin if(four_bit_hash == 0) next_state = 1035; else  next_state = 2000;  end 
1035: begin if(four_bit_hash == 0) next_state = 1036; else  next_state = 2000;  end 
1036: begin if(four_bit_hash == 0) next_state = 1037; else  next_state = 2000;  end 
1037: begin if(four_bit_hash == 0) next_state = 1038; else  next_state = 2000;  end 
1038: begin if(four_bit_hash == 0) next_state = 1039; else  next_state = 2000;  end 
1039: begin if(four_bit_hash == 0) next_state = 1040; else  next_state = 2000;  end 
1040: begin if(four_bit_hash == 0) next_state = 1041; else  next_state = 2000;  end 
1041: begin if(four_bit_hash == 0) next_state = 1042; else  next_state = 2000;  end 
1042: begin if(four_bit_hash == 0) next_state = 1043; else  next_state = 2000;  end 
1043: begin if(four_bit_hash == 0) next_state = 1044; else  next_state = 2000;  end 
1044: begin if(four_bit_hash == 0) next_state = 1045; else  next_state = 2000;  end 
1045: begin if(four_bit_hash == 0) next_state = 1046; else  next_state = 2000;  end 
1046: begin if(four_bit_hash == 0) next_state = 1047; else  next_state = 2000;  end 
1047: begin if(four_bit_hash == 0) next_state = 1048; else  next_state = 2000;  end 
1048: begin if(four_bit_hash == 0) next_state = 1049; else  next_state = 2000;  end 
1049: begin if(four_bit_hash == 0) next_state = 1050; else  next_state = 2000;  end 
1050: begin if(four_bit_hash == 0) next_state = 1051; else  next_state = 2000;  end 
1051: begin if(four_bit_hash == 0) next_state = 1052; else  next_state = 2000;  end 
1052: begin if(four_bit_hash == 0) next_state = 1053; else  next_state = 2000;  end 
1053: begin if(four_bit_hash == 0) next_state = 1054; else  next_state = 2000;  end 
1054: begin if(four_bit_hash == 0) next_state = 1055; else  next_state = 2000;  end 
1055: begin if(four_bit_hash == 0) next_state = 1056; else  next_state = 2000;  end 
1056: begin if(four_bit_hash == 0) next_state = 1057; else  next_state = 2000;  end 
1057: begin if(four_bit_hash == 0) next_state = 1058; else  next_state = 2000;  end 
1058: begin if(four_bit_hash == 0) next_state = 1059; else  next_state = 2000;  end 
1059: begin if(four_bit_hash == 0) next_state = 1060; else  next_state = 2000;  end 
1060: begin if(four_bit_hash == 0) next_state = 1061; else  next_state = 2000;  end 
1061: begin if(four_bit_hash == 0) next_state = 1062; else  next_state = 2000;  end 
1062: begin if(four_bit_hash == 0) next_state = 1063; else  next_state = 2000;  end 
1063: begin if(four_bit_hash == 0) next_state = 1064; else  next_state = 2000;  end 
1064: begin if(four_bit_hash == 0) next_state = 1065; else  next_state = 2000;  end 
1065: begin if(four_bit_hash == 0) next_state = 1066; else  next_state = 2000;  end 
1066: begin if(four_bit_hash == 0) next_state = 1067; else  next_state = 2000;  end 
1067: begin if(four_bit_hash == 0) next_state = 1068; else  next_state = 2000;  end 
1068: begin if(four_bit_hash == 0) next_state = 1069; else  next_state = 2000;  end 
1069: begin if(four_bit_hash == 0) next_state = 1070; else  next_state = 2000;  end 
1070: begin if(four_bit_hash == 0) next_state = 1071; else  next_state = 2000;  end 
1071: begin if(four_bit_hash == 0) next_state = 1072; else  next_state = 2000;  end 
1072: begin if(four_bit_hash == 0) next_state = 1073; else  next_state = 2000;  end 
1073: begin if(four_bit_hash == 0) next_state = 1074; else  next_state = 2000;  end 
1074: begin if(four_bit_hash == 0) next_state = 1075; else  next_state = 2000;  end 
1075: begin if(four_bit_hash == 0) next_state = 1076; else  next_state = 2000;  end 
1076: begin if(four_bit_hash == 0) next_state = 1077; else  next_state = 2000;  end 
1077: begin if(four_bit_hash == 0) next_state = 1078; else  next_state = 2000;  end 
1078: begin if(four_bit_hash == 0) next_state = 1079; else  next_state = 2000;  end 
1079: begin if(four_bit_hash == 0) next_state = 1080; else  next_state = 2000;  end 
1080: begin if(four_bit_hash == 0) next_state = 1081; else  next_state = 2000;  end 
1081: begin if(four_bit_hash == 0) next_state = 1082; else  next_state = 2000;  end 
1082: begin if(four_bit_hash == 0) next_state = 1083; else  next_state = 2000;  end 
1083: begin if(four_bit_hash == 0) next_state = 1084; else  next_state = 2000;  end 
1084: begin if(four_bit_hash == 0) next_state = 1085; else  next_state = 2000;  end 
1085: begin if(four_bit_hash == 0) next_state = 1086; else  next_state = 2000;  end 
1086: begin if(four_bit_hash == 0) next_state = 1087; else  next_state = 2000;  end 
1087: begin if(four_bit_hash == 0) next_state = 1088; else  next_state = 2000;  end 
1088: begin if(four_bit_hash == 0) next_state = 1089; else  next_state = 2000;  end 
1089: begin if(four_bit_hash == 0) next_state = 1090; else  next_state = 2000;  end 
1090: begin if(four_bit_hash == 0) next_state = 1091; else  next_state = 2000;  end 
1091: begin if(four_bit_hash == 0) next_state = 1092; else  next_state = 2000;  end 
1092: begin if(four_bit_hash == 0) next_state = 1093; else  next_state = 2000;  end 
1093: begin if(four_bit_hash == 0) next_state = 1094; else  next_state = 2000;  end 
1094: begin if(four_bit_hash == 0) next_state = 1095; else  next_state = 2000;  end 
1095: begin if(four_bit_hash == 0) next_state = 1096; else  next_state = 2000;  end 
1096: begin if(four_bit_hash == 0) next_state = 1097; else  next_state = 2000;  end 
1097: begin if(four_bit_hash == 0) next_state = 1098; else  next_state = 2000;  end 
1098: begin if(four_bit_hash == 0) next_state = 1099; else  next_state = 2000;  end 
1099: begin if(four_bit_hash == 0) next_state = 1100; else  next_state = 2000;  end 
1100: begin if(four_bit_hash == 0) next_state = 1101; else  next_state = 2000;  end 
1101: begin if(four_bit_hash == 0) next_state = 1102; else  next_state = 2000;  end 
1102: begin if(four_bit_hash == 0) next_state = 1103; else  next_state = 2000;  end 
1103: begin if(four_bit_hash == 0) next_state = 1104; else  next_state = 2000;  end 
1104: begin if(four_bit_hash == 0) next_state = 1105; else  next_state = 2000;  end 
1105: begin if(four_bit_hash == 0) next_state = 1106; else  next_state = 2000;  end 
1106: begin if(four_bit_hash == 0) next_state = 1107; else  next_state = 2000;  end 
1107: begin if(four_bit_hash == 0) next_state = 1108; else  next_state = 2000;  end 
1108: begin if(four_bit_hash == 0) next_state = 1109; else  next_state = 2000;  end 
1109: begin if(four_bit_hash == 0) next_state = 1110; else  next_state = 2000;  end 
1110: begin if(four_bit_hash == 0) next_state = 1111; else  next_state = 2000;  end 
1111: begin if(four_bit_hash == 0) next_state = 1112; else  next_state = 2000;  end 
1112: begin if(four_bit_hash == 0) next_state = 1113; else  next_state = 2000;  end 
1113: begin if(four_bit_hash == 0) next_state = 1114; else  next_state = 2000;  end 
1114: begin if(four_bit_hash == 0) next_state = 1115; else  next_state = 2000;  end 
1115: begin if(four_bit_hash == 0) next_state = 1116; else  next_state = 2000;  end 
1116: begin if(four_bit_hash == 0) next_state = 1117; else  next_state = 2000;  end 
1117: begin if(four_bit_hash == 0) next_state = 1118; else  next_state = 2000;  end 
1118: begin if(four_bit_hash == 0) next_state = 1119; else  next_state = 2000;  end 
1119: begin if(four_bit_hash == 0) next_state = 1120; else  next_state = 2000;  end 
1120: begin if(four_bit_hash == 0) next_state = 1121; else  next_state = 2000;  end 
1121: begin if(four_bit_hash == 0) next_state = 1122; else  next_state = 2000;  end 
1122: begin if(four_bit_hash == 0) next_state = 1123; else  next_state = 2000;  end 
1123: begin if(four_bit_hash == 0) next_state = 1124; else  next_state = 2000;  end 
1124: begin if(four_bit_hash == 0) next_state = 1125; else  next_state = 2000;  end 
1125: begin if(four_bit_hash == 0) next_state = 1126; else  next_state = 2000;  end 
1126: begin if(four_bit_hash == 0) next_state = 1127; else  next_state = 2000;  end 
1127: begin if(four_bit_hash == 0) next_state = 1128; else  next_state = 2000;  end 
1128: begin if(four_bit_hash == 0) next_state = 1129; else  next_state = 2000;  end 
1129: begin if(four_bit_hash == 0) next_state = 1130; else  next_state = 2000;  end 
1130: begin if(four_bit_hash == 0) next_state = 1131; else  next_state = 2000;  end 
1131: begin if(four_bit_hash == 0) next_state = 1132; else  next_state = 2000;  end 
1132: begin if(four_bit_hash == 0) next_state = 1133; else  next_state = 2000;  end 
1133: begin if(four_bit_hash == 0) next_state = 1134; else  next_state = 2000;  end 
1134: begin if(four_bit_hash == 0) next_state = 1135; else  next_state = 2000;  end 
1135: begin if(four_bit_hash == 0) next_state = 1136; else  next_state = 2000;  end 
1136: begin if(four_bit_hash == 0) next_state = 1137; else  next_state = 2000;  end 
1137: begin if(four_bit_hash == 0) next_state = 1138; else  next_state = 2000;  end 
1138: begin if(four_bit_hash == 0) next_state = 1139; else  next_state = 2000;  end 
1139: begin if(four_bit_hash == 0) next_state = 1140; else  next_state = 2000;  end 
1140: begin if(four_bit_hash == 0) next_state = 1141; else  next_state = 2000;  end 
1141: begin if(four_bit_hash == 0) next_state = 1142; else  next_state = 2000;  end 
1142: begin if(four_bit_hash == 0) next_state = 1143; else  next_state = 2000;  end 
1143: begin if(four_bit_hash == 0) next_state = 1144; else  next_state = 2000;  end 
1144: begin if(four_bit_hash == 0) next_state = 1145; else  next_state = 2000;  end 
1145: begin if(four_bit_hash == 0) next_state = 1146; else  next_state = 2000;  end 
1146: begin if(four_bit_hash == 0) next_state = 1147; else  next_state = 2000;  end 
1147: begin if(four_bit_hash == 0) next_state = 1148; else  next_state = 2000;  end 
1148: begin if(four_bit_hash == 0) next_state = 1149; else  next_state = 2000;  end 
1149: begin if(four_bit_hash == 0) next_state = 1150; else  next_state = 2000;  end 
1150: begin if(four_bit_hash == 0) next_state = 1151; else  next_state = 2000;  end 
1151: begin if(four_bit_hash == 0) next_state = 1152; else  next_state = 2000;  end 
1152: begin if(four_bit_hash == 0) next_state = 1153; else  next_state = 2000;  end 
1153: begin if(four_bit_hash == 0) next_state = 1154; else  next_state = 2000;  end 
1154: begin if(four_bit_hash == 0) next_state = 1155; else  next_state = 2000;  end 
1155: begin if(four_bit_hash == 0) next_state = 1156; else  next_state = 2000;  end 
1156: begin if(four_bit_hash == 0) next_state = 1157; else  next_state = 2000;  end 
1157: begin if(four_bit_hash == 0) next_state = 1158; else  next_state = 2000;  end 
1158: begin if(four_bit_hash == 0) next_state = 1159; else  next_state = 2000;  end 
1159: begin if(four_bit_hash == 0) next_state = 1160; else  next_state = 2000;  end 
1160: begin if(four_bit_hash == 0) next_state = 1161; else  next_state = 2000;  end 
1161: begin if(four_bit_hash == 0) next_state = 1162; else  next_state = 2000;  end 
1162: begin if(four_bit_hash == 0) next_state = 1163; else  next_state = 2000;  end 
1163: begin if(four_bit_hash == 0) next_state = 1164; else  next_state = 2000;  end 
1164: begin if(four_bit_hash == 0) next_state = 1165; else  next_state = 2000;  end 
1165: begin if(four_bit_hash == 0) next_state = 1166; else  next_state = 2000;  end 
1166: begin if(four_bit_hash == 0) next_state = 1167; else  next_state = 2000;  end 
1167: begin if(four_bit_hash == 0) next_state = 1168; else  next_state = 2000;  end 
1168: begin if(four_bit_hash == 0) next_state = 1169; else  next_state = 2000;  end 
1169: begin if(four_bit_hash == 0) next_state = 1170; else  next_state = 2000;  end 
1170: begin if(four_bit_hash == 0) next_state = 1171; else  next_state = 2000;  end 
1171: begin if(four_bit_hash == 0) next_state = 1172; else  next_state = 2000;  end 
1172: begin if(four_bit_hash == 0) next_state = 1173; else  next_state = 2000;  end 
1173: begin if(four_bit_hash == 0) next_state = 1174; else  next_state = 2000;  end 
1174: begin if(four_bit_hash == 0) next_state = 1175; else  next_state = 2000;  end 
1175: begin if(four_bit_hash == 0) next_state = 1176; else  next_state = 2000;  end 
1176: begin if(four_bit_hash == 0) next_state = 1177; else  next_state = 2000;  end 
1177: begin if(four_bit_hash == 0) next_state = 1178; else  next_state = 2000;  end 
1178: begin if(four_bit_hash == 0) next_state = 1179; else  next_state = 2000;  end 
1179: begin if(four_bit_hash == 0) next_state = 1180; else  next_state = 2000;  end 
1180: begin if(four_bit_hash == 0) next_state = 1181; else  next_state = 2000;  end 
1181: begin if(four_bit_hash == 0) next_state = 1182; else  next_state = 2000;  end 
1182: begin if(four_bit_hash == 0) next_state = 1183; else  next_state = 2000;  end 
1183: begin if(four_bit_hash == 0) next_state = 1184; else  next_state = 2000;  end 
1184: begin if(four_bit_hash == 0) next_state = 1185; else  next_state = 2000;  end 
1185: begin if(four_bit_hash == 0) next_state = 1186; else  next_state = 2000;  end 
1186: begin if(four_bit_hash == 0) next_state = 1187; else  next_state = 2000;  end 
1187: begin if(four_bit_hash == 0) next_state = 1188; else  next_state = 2000;  end 
1188: begin if(four_bit_hash == 0) next_state = 1189; else  next_state = 2000;  end 
1189: begin if(four_bit_hash == 0) next_state = 1190; else  next_state = 2000;  end 
1190: begin if(four_bit_hash == 0) next_state = 1191; else  next_state = 2000;  end 
1191: begin if(four_bit_hash == 0) next_state = 1192; else  next_state = 2000;  end 
1192: begin if(four_bit_hash == 0) next_state = 1193; else  next_state = 2000;  end 
1193: begin if(four_bit_hash == 0) next_state = 1194; else  next_state = 2000;  end 
1194: begin if(four_bit_hash == 0) next_state = 1195; else  next_state = 2000;  end 
1195: begin if(four_bit_hash == 0) next_state = 1196; else  next_state = 2000;  end 
1196: begin if(four_bit_hash == 0) next_state = 1197; else  next_state = 2000;  end 
1197: begin if(four_bit_hash == 0) next_state = 1198; else  next_state = 2000;  end 
1198: begin if(four_bit_hash == 0) next_state = 1199; else  next_state = 2000;  end 
1199: begin if(four_bit_hash == 0) next_state = 1200; else  next_state = 2000;  end 
1200: begin if(four_bit_hash == 0) next_state = 1201; else  next_state = 2000;  end 
1201: begin if(four_bit_hash == 0) next_state = 1202; else  next_state = 2000;  end 
1202: begin if(four_bit_hash == 0) next_state = 1203; else  next_state = 2000;  end 
1203: begin if(four_bit_hash == 0) next_state = 1204; else  next_state = 2000;  end 
1204: begin if(four_bit_hash == 0) next_state = 1205; else  next_state = 2000;  end 
1205: begin if(four_bit_hash == 0) next_state = 1206; else  next_state = 2000;  end 
1206: begin if(four_bit_hash == 0) next_state = 1207; else  next_state = 2000;  end 
1207: begin if(four_bit_hash == 0) next_state = 1208; else  next_state = 2000;  end 
1208: begin if(four_bit_hash == 0) next_state = 1209; else  next_state = 2000;  end 
1209: begin if(four_bit_hash == 0) next_state = 1210; else  next_state = 2000;  end 
1210: begin if(four_bit_hash == 0) next_state = 1211; else  next_state = 2000;  end 
1211: begin if(four_bit_hash == 0) next_state = 1212; else  next_state = 2000;  end 
1212: begin if(four_bit_hash == 0) next_state = 1213; else  next_state = 2000;  end 
1213: begin if(four_bit_hash == 0) next_state = 1214; else  next_state = 2000;  end 
1214: begin if(four_bit_hash == 0) next_state = 1215; else  next_state = 2000;  end 
1215: begin if(four_bit_hash == 0) next_state = 1216; else  next_state = 2000;  end 
1216: begin if(four_bit_hash == 0) next_state = 1217; else  next_state = 2000;  end 
1217: begin if(four_bit_hash == 0) next_state = 1218; else  next_state = 2000;  end 
1218: begin if(four_bit_hash == 0) next_state = 1219; else  next_state = 2000;  end 
1219: begin if(four_bit_hash == 0) next_state = 1220; else  next_state = 2000;  end 
1220: begin if(four_bit_hash == 0) next_state = 1221; else  next_state = 2000;  end 
1221: begin if(four_bit_hash == 0) next_state = 1222; else  next_state = 2000;  end 
1222: begin if(four_bit_hash == 0) next_state = 1223; else  next_state = 2000;  end 
1223: begin if(four_bit_hash == 0) next_state = 1224; else  next_state = 2000;  end 
1224: begin if(four_bit_hash == 0) next_state = 1225; else  next_state = 2000;  end 
1225: begin if(four_bit_hash == 0) next_state = 1226; else  next_state = 2000;  end 
1226: begin if(four_bit_hash == 0) next_state = 1227; else  next_state = 2000;  end 
1227: begin if(four_bit_hash == 0) next_state = 1228; else  next_state = 2000;  end 
1228: begin if(four_bit_hash == 0) next_state = 1229; else  next_state = 2000;  end 
1229: begin if(four_bit_hash == 0) next_state = 1230; else  next_state = 2000;  end 
1230: begin if(four_bit_hash == 0) next_state = 1231; else  next_state = 2000;  end 
1231: begin if(four_bit_hash == 0) next_state = 1232; else  next_state = 2000;  end 
1232: begin if(four_bit_hash == 0) next_state = 1233; else  next_state = 2000;  end 
1233: begin if(four_bit_hash == 0) next_state = 1234; else  next_state = 2000;  end 
1234: begin if(four_bit_hash == 0) next_state = 1235; else  next_state = 2000;  end 
1235: begin if(four_bit_hash == 0) next_state = 1236; else  next_state = 2000;  end 
1236: begin if(four_bit_hash == 0) next_state = 1237; else  next_state = 2000;  end 
1237: begin if(four_bit_hash == 0) next_state = 1238; else  next_state = 2000;  end 
1238: begin if(four_bit_hash == 0) next_state = 1239; else  next_state = 2000;  end 
1239: begin if(four_bit_hash == 0) next_state = 1240; else  next_state = 2000;  end 
1240: begin if(four_bit_hash == 0) next_state = 1241; else  next_state = 2000;  end 
1241: begin if(four_bit_hash == 0) next_state = 1242; else  next_state = 2000;  end 
1242: begin if(four_bit_hash == 0) next_state = 1243; else  next_state = 2000;  end 
1243: begin if(four_bit_hash == 0) next_state = 1244; else  next_state = 2000;  end 
1244: begin if(four_bit_hash == 0) next_state = 1245; else  next_state = 2000;  end 
1245: begin if(four_bit_hash == 0) next_state = 1246; else  next_state = 2000;  end 
1246: begin if(four_bit_hash == 0) next_state = 1247; else  next_state = 2000;  end 
1247: begin if(four_bit_hash == 0) next_state = 1248; else  next_state = 2000;  end 
1248: begin if(four_bit_hash == 0) next_state = 1249; else  next_state = 2000;  end 
1249: begin if(four_bit_hash == 0) next_state = 1250; else  next_state = 2000;  end 
1250: begin if(four_bit_hash == 0) next_state = 1251; else  next_state = 2000;  end 
1251: begin if(four_bit_hash == 0) next_state = 1252; else  next_state = 2000;  end 
1252: begin if(four_bit_hash == 0) next_state = 1253; else  next_state = 2000;  end 
1253: begin if(four_bit_hash == 0) next_state = 1254; else  next_state = 2000;  end 
1254: begin if(four_bit_hash == 0) next_state = 1255; else  next_state = 2000;  end 
1255: begin if(four_bit_hash == 0) next_state = 1256; else  next_state = 2000;  end 
1256: begin if(four_bit_hash == 0) next_state = 1257; else  next_state = 2000;  end 
1257: begin if(four_bit_hash == 0) next_state = 1258; else  next_state = 2000;  end 
1258: begin if(four_bit_hash == 0) next_state = 1259; else  next_state = 2000;  end 
1259: begin if(four_bit_hash == 0) next_state = 1260; else  next_state = 2000;  end 
1260: begin if(four_bit_hash == 0) next_state = 1261; else  next_state = 2000;  end 
1261: begin if(four_bit_hash == 0) next_state = 1262; else  next_state = 2000;  end 
1262: begin if(four_bit_hash == 0) next_state = 1263; else  next_state = 2000;  end 
1263: begin if(four_bit_hash == 0) next_state = 1264; else  next_state = 2000;  end 
1264: begin if(four_bit_hash == 0) next_state = 1265; else  next_state = 2000;  end 
1265: begin if(four_bit_hash == 0) next_state = 1266; else  next_state = 2000;  end 
1266: begin if(four_bit_hash == 0) next_state = 1267; else  next_state = 2000;  end 
1267: begin if(four_bit_hash == 0) next_state = 1268; else  next_state = 2000;  end 
1268: begin if(four_bit_hash == 0) next_state = 1269; else  next_state = 2000;  end 
1269: begin if(four_bit_hash == 0) next_state = 1270; else  next_state = 2000;  end 
1270: begin if(four_bit_hash == 0) next_state = 1271; else  next_state = 2000;  end 
1271: begin if(four_bit_hash == 0) next_state = 1272; else  next_state = 2000;  end 
1272: begin if(four_bit_hash == 0) next_state = 1273; else  next_state = 2000;  end 
1273: begin if(four_bit_hash == 0) next_state = 1274; else  next_state = 2000;  end 
1274: begin if(four_bit_hash == 0) next_state = 1275; else  next_state = 2000;  end 
1275: begin if(four_bit_hash == 0) next_state = 1276; else  next_state = 2000;  end 
1276: begin if(four_bit_hash == 0) next_state = 1277; else  next_state = 2000;  end 
1277: begin if(four_bit_hash == 0) next_state = 1278; else  next_state = 2000;  end 
1278: begin if(four_bit_hash == 0) next_state = 1279; else  next_state = 2000;  end 
1279: begin if(four_bit_hash == 0) next_state = 1280; else  next_state = 2000;  end 
1280: begin if(four_bit_hash == 0) next_state = 1281; else  next_state = 2000;  end 
1281: begin if(four_bit_hash == 0) next_state = 1282; else  next_state = 2000;  end 
1282: begin if(four_bit_hash == 0) next_state = 1283; else  next_state = 2000;  end 
1283: begin if(four_bit_hash == 0) next_state = 1284; else  next_state = 2000;  end 
1284: begin if(four_bit_hash == 0) next_state = 1285; else  next_state = 2000;  end 
1285: begin if(four_bit_hash == 0) next_state = 1286; else  next_state = 2000;  end 
1286: begin if(four_bit_hash == 0) next_state = 1287; else  next_state = 2000;  end 
1287: begin if(four_bit_hash == 0) next_state = 1288; else  next_state = 2000;  end 
1288: begin if(four_bit_hash == 0) next_state = 1289; else  next_state = 2000;  end 
1289: begin if(four_bit_hash == 0) next_state = 1290; else  next_state = 2000;  end 
1290: begin if(four_bit_hash == 0) next_state = 1291; else  next_state = 2000;  end 
1291: begin if(four_bit_hash == 0) next_state = 1292; else  next_state = 2000;  end 
1292: begin if(four_bit_hash == 0) next_state = 1293; else  next_state = 2000;  end 
1293: begin if(four_bit_hash == 0) next_state = 1294; else  next_state = 2000;  end 
1294: begin if(four_bit_hash == 0) next_state = 1295; else  next_state = 2000;  end 
1295: begin if(four_bit_hash == 0) next_state = 1296; else  next_state = 2000;  end 
1296: begin if(four_bit_hash == 0) next_state = 1297; else  next_state = 2000;  end 
1297: begin if(four_bit_hash == 0) next_state = 1298; else  next_state = 2000;  end 
1298: begin if(four_bit_hash == 0) next_state = 1299; else  next_state = 2000;  end 
1299: begin if(four_bit_hash == 0) next_state = 1300; else  next_state = 2000;  end 
1300: begin if(four_bit_hash == 0) next_state = 1301; else  next_state = 2000;  end 
1301: begin if(four_bit_hash == 0) next_state = 1302; else  next_state = 2000;  end 
1302: begin if(four_bit_hash == 0) next_state = 1303; else  next_state = 2000;  end 
1303: begin if(four_bit_hash == 0) next_state = 1304; else  next_state = 2000;  end 
1304: begin if(four_bit_hash == 0) next_state = 1305; else  next_state = 2000;  end 
1305: begin if(four_bit_hash == 0) next_state = 1306; else  next_state = 2000;  end 
1306: begin if(four_bit_hash == 0) next_state = 1307; else  next_state = 2000;  end 
1307: begin if(four_bit_hash == 0) next_state = 1308; else  next_state = 2000;  end 
1308: begin if(four_bit_hash == 0) next_state = 1309; else  next_state = 2000;  end 
1309: begin if(four_bit_hash == 0) next_state = 1310; else  next_state = 2000;  end 
1310: begin if(four_bit_hash == 0) next_state = 1311; else  next_state = 2000;  end 
1311: begin if(four_bit_hash == 0) next_state = 1312; else  next_state = 2000;  end 
1312: begin if(four_bit_hash == 0) next_state = 1313; else  next_state = 2000;  end 
1313: begin if(four_bit_hash == 0) next_state = 1314; else  next_state = 2000;  end 
1314: begin if(four_bit_hash == 0) next_state = 1315; else  next_state = 2000;  end 
1315: begin if(four_bit_hash == 0) next_state = 1316; else  next_state = 2000;  end 
1316: begin if(four_bit_hash == 0) next_state = 1317; else  next_state = 2000;  end 
1317: begin if(four_bit_hash == 0) next_state = 1318; else  next_state = 2000;  end 
1318: begin if(four_bit_hash == 0) next_state = 1319; else  next_state = 2000;  end 
1319: begin if(four_bit_hash == 0) next_state = 1320; else  next_state = 2000;  end 
1320: begin if(four_bit_hash == 0) next_state = 1321; else  next_state = 2000;  end 
1321: begin if(four_bit_hash == 0) next_state = 1322; else  next_state = 2000;  end 
1322: begin if(four_bit_hash == 0) next_state = 1323; else  next_state = 2000;  end 
1323: begin if(four_bit_hash == 0) next_state = 1324; else  next_state = 2000;  end 
1324: begin if(four_bit_hash == 0) next_state = 1325; else  next_state = 2000;  end 
1325: begin if(four_bit_hash == 0) next_state = 1326; else  next_state = 2000;  end 
1326: begin if(four_bit_hash == 0) next_state = 1327; else  next_state = 2000;  end 
1327: begin if(four_bit_hash == 0) next_state = 1328; else  next_state = 2000;  end 
1328: begin if(four_bit_hash == 0) next_state = 1329; else  next_state = 2000;  end 
1329: begin if(four_bit_hash == 0) next_state = 1330; else  next_state = 2000;  end 
1330: begin if(four_bit_hash == 0) next_state = 1331; else  next_state = 2000;  end 
1331: begin if(four_bit_hash == 0) next_state = 1332; else  next_state = 2000;  end 
1332: begin if(four_bit_hash == 0) next_state = 1333; else  next_state = 2000;  end 
1333: begin if(four_bit_hash == 0) next_state = 1334; else  next_state = 2000;  end 
1334: begin if(four_bit_hash == 0) next_state = 1335; else  next_state = 2000;  end 
1335: begin if(four_bit_hash == 0) next_state = 1336; else  next_state = 2000;  end 
1336: begin if(four_bit_hash == 0) next_state = 1337; else  next_state = 2000;  end 
1337: begin if(four_bit_hash == 0) next_state = 1338; else  next_state = 2000;  end 
1338: begin if(four_bit_hash == 0) next_state = 1339; else  next_state = 2000;  end 
1339: begin if(four_bit_hash == 0) next_state = 1340; else  next_state = 2000;  end 
1340: begin if(four_bit_hash == 0) next_state = 1341; else  next_state = 2000;  end 
1341: begin if(four_bit_hash == 0) next_state = 1342; else  next_state = 2000;  end 
1342: begin if(four_bit_hash == 0) next_state = 1343; else  next_state = 2000;  end 
1343: begin if(four_bit_hash == 0) next_state = 1344; else  next_state = 2000;  end 
1344: begin if(four_bit_hash == 0) next_state = 1345; else  next_state = 2000;  end 
1345: begin if(four_bit_hash == 0) next_state = 1346; else  next_state = 2000;  end 
1346: begin if(four_bit_hash == 0) next_state = 1347; else  next_state = 2000;  end 
1347: begin if(four_bit_hash == 0) next_state = 1348; else  next_state = 2000;  end 
1348: begin if(four_bit_hash == 0) next_state = 1349; else  next_state = 2000;  end 
1349: begin if(four_bit_hash == 0) next_state = 1350; else  next_state = 2000;  end 
1350: begin if(four_bit_hash == 0) next_state = 1351; else  next_state = 2000;  end 
1351: begin if(four_bit_hash == 0) next_state = 1352; else  next_state = 2000;  end 
1352: begin if(four_bit_hash == 0) next_state = 1353; else  next_state = 2000;  end 
1353: begin if(four_bit_hash == 0) next_state = 1354; else  next_state = 2000;  end 
1354: begin if(four_bit_hash == 0) next_state = 1355; else  next_state = 2000;  end 
1355: begin if(four_bit_hash == 0) next_state = 1356; else  next_state = 2000;  end 
1356: begin if(four_bit_hash == 0) next_state = 1357; else  next_state = 2000;  end 
1357: begin if(four_bit_hash == 0) next_state = 1358; else  next_state = 2000;  end 
1358: begin if(four_bit_hash == 0) next_state = 1359; else  next_state = 2000;  end 
1359: begin if(four_bit_hash == 0) next_state = 1360; else  next_state = 2000;  end 
1360: begin if(four_bit_hash == 0) next_state = 1361; else  next_state = 2000;  end 
1361: begin if(four_bit_hash == 0) next_state = 1362; else  next_state = 2000;  end 
1362: begin if(four_bit_hash == 0) next_state = 1363; else  next_state = 2000;  end 
1363: begin if(four_bit_hash == 0) next_state = 1364; else  next_state = 2000;  end 
1364: begin if(four_bit_hash == 0) next_state = 1365; else  next_state = 2000;  end 
1365: begin if(four_bit_hash == 0) next_state = 1366; else  next_state = 2000;  end 
1366: begin if(four_bit_hash == 0) next_state = 1367; else  next_state = 2000;  end 
1367: begin if(four_bit_hash == 0) next_state = 1368; else  next_state = 2000;  end 
1368: begin if(four_bit_hash == 0) next_state = 1369; else  next_state = 2000;  end 
1369: begin if(four_bit_hash == 0) next_state = 1370; else  next_state = 2000;  end 
1370: begin if(four_bit_hash == 0) next_state = 1371; else  next_state = 2000;  end 
1371: begin if(four_bit_hash == 0) next_state = 1372; else  next_state = 2000;  end 
1372: begin if(four_bit_hash == 0) next_state = 1373; else  next_state = 2000;  end 
1373: begin if(four_bit_hash == 0) next_state = 1374; else  next_state = 2000;  end 
1374: begin if(four_bit_hash == 0) next_state = 1375; else  next_state = 2000;  end 
1375: begin if(four_bit_hash == 0) next_state = 1376; else  next_state = 2000;  end 
1376: begin if(four_bit_hash == 0) next_state = 1377; else  next_state = 2000;  end 
1377: begin if(four_bit_hash == 0) next_state = 1378; else  next_state = 2000;  end 
1378: begin if(four_bit_hash == 0) next_state = 1379; else  next_state = 2000;  end 
1379: begin if(four_bit_hash == 0) next_state = 1380; else  next_state = 2000;  end 
1380: begin if(four_bit_hash == 0) next_state = 1381; else  next_state = 2000;  end 
1381: begin if(four_bit_hash == 0) next_state = 1382; else  next_state = 2000;  end 
1382: begin if(four_bit_hash == 0) next_state = 1383; else  next_state = 2000;  end 
1383: begin if(four_bit_hash == 0) next_state = 1384; else  next_state = 2000;  end 
1384: begin if(four_bit_hash == 0) next_state = 1385; else  next_state = 2000;  end 
1385: begin if(four_bit_hash == 0) next_state = 1386; else  next_state = 2000;  end 
1386: begin if(four_bit_hash == 0) next_state = 1387; else  next_state = 2000;  end 
1387: begin if(four_bit_hash == 0) next_state = 1388; else  next_state = 2000;  end 
1388: begin if(four_bit_hash == 0) next_state = 1389; else  next_state = 2000;  end 
1389: begin if(four_bit_hash == 0) next_state = 1390; else  next_state = 2000;  end 
1390: begin if(four_bit_hash == 0) next_state = 1391; else  next_state = 2000;  end 
1391: begin if(four_bit_hash == 0) next_state = 1392; else  next_state = 2000;  end 
1392: begin if(four_bit_hash == 0) next_state = 1393; else  next_state = 2000;  end 
1393: begin if(four_bit_hash == 0) next_state = 1394; else  next_state = 2000;  end 
1394: begin if(four_bit_hash == 0) next_state = 1395; else  next_state = 2000;  end 
1395: begin if(four_bit_hash == 0) next_state = 1396; else  next_state = 2000;  end 
1396: begin if(four_bit_hash == 0) next_state = 1397; else  next_state = 2000;  end 
1397: begin if(four_bit_hash == 0) next_state = 1398; else  next_state = 2000;  end 
1398: begin if(four_bit_hash == 0) next_state = 1399; else  next_state = 2000;  end 
1399: begin if(four_bit_hash == 0) next_state = 1400; else  next_state = 2000;  end 
1400: begin if(four_bit_hash == 0) next_state = 1401; else  next_state = 2000;  end 
1401: begin if(four_bit_hash == 0) next_state = 1402; else  next_state = 2000;  end 
1402: begin if(four_bit_hash == 0) next_state = 1403; else  next_state = 2000;  end 
1403: begin if(four_bit_hash == 0) next_state = 1404; else  next_state = 2000;  end 
1404: begin if(four_bit_hash == 0) next_state = 1405; else  next_state = 2000;  end 
1405: begin if(four_bit_hash == 0) next_state = 1406; else  next_state = 2000;  end 
1406: begin if(four_bit_hash == 0) next_state = 1407; else  next_state = 2000;  end 
1407: begin if(four_bit_hash == 0) next_state = 1408; else  next_state = 2000;  end 
1408: begin if(four_bit_hash == 0) next_state = 1409; else  next_state = 2000;  end 
1409: begin if(four_bit_hash == 0) next_state = 1410; else  next_state = 2000;  end 
1410: begin if(four_bit_hash == 0) next_state = 1411; else  next_state = 2000;  end 
1411: begin if(four_bit_hash == 0) next_state = 1412; else  next_state = 2000;  end 
1412: begin if(four_bit_hash == 0) next_state = 1413; else  next_state = 2000;  end 
1413: begin if(four_bit_hash == 0) next_state = 1414; else  next_state = 2000;  end 
1414: begin if(four_bit_hash == 0) next_state = 1415; else  next_state = 2000;  end 
1415: begin if(four_bit_hash == 0) next_state = 1416; else  next_state = 2000;  end 
1416: begin if(four_bit_hash == 0) next_state = 1417; else  next_state = 2000;  end 
1417: begin if(four_bit_hash == 0) next_state = 1418; else  next_state = 2000;  end 
1418: begin if(four_bit_hash == 0) next_state = 1419; else  next_state = 2000;  end 
1419: begin if(four_bit_hash == 0) next_state = 1420; else  next_state = 2000;  end 
1420: begin if(four_bit_hash == 0) next_state = 1421; else  next_state = 2000;  end 
1421: begin if(four_bit_hash == 0) next_state = 1422; else  next_state = 2000;  end 
1422: begin if(four_bit_hash == 0) next_state = 1423; else  next_state = 2000;  end 
1423: begin if(four_bit_hash == 0) next_state = 1424; else  next_state = 2000;  end 
1424: begin if(four_bit_hash == 0) next_state = 1425; else  next_state = 2000;  end 
1425: begin if(four_bit_hash == 0) next_state = 1426; else  next_state = 2000;  end 
1426: begin if(four_bit_hash == 0) next_state = 1427; else  next_state = 2000;  end 
1427: begin if(four_bit_hash == 0) next_state = 1428; else  next_state = 2000;  end 
1428: begin if(four_bit_hash == 0) next_state = 1429; else  next_state = 2000;  end 
1429: begin if(four_bit_hash == 0) next_state = 1430; else  next_state = 2000;  end 
1430: begin if(four_bit_hash == 0) next_state = 1431; else  next_state = 2000;  end 
1431: begin if(four_bit_hash == 0) next_state = 1432; else  next_state = 2000;  end 
1432: begin if(four_bit_hash == 0) next_state = 1433; else  next_state = 2000;  end 
1433: begin if(four_bit_hash == 0) next_state = 1434; else  next_state = 2000;  end 
1434: begin if(four_bit_hash == 0) next_state = 1435; else  next_state = 2000;  end 
1435: begin if(four_bit_hash == 0) next_state = 1436; else  next_state = 2000;  end 
1436: begin if(four_bit_hash == 0) next_state = 1437; else  next_state = 2000;  end 
1437: begin if(four_bit_hash == 0) next_state = 1438; else  next_state = 2000;  end 
1438: begin if(four_bit_hash == 0) next_state = 1439; else  next_state = 2000;  end 
1439: begin if(four_bit_hash == 0) next_state = 1440; else  next_state = 2000;  end 
1440: begin if(four_bit_hash == 0) next_state = 1441; else  next_state = 2000;  end 
1441: begin if(four_bit_hash == 0) next_state = 1442; else  next_state = 2000;  end 
1442: begin if(four_bit_hash == 0) next_state = 1443; else  next_state = 2000;  end 
1443: begin if(four_bit_hash == 0) next_state = 1444; else  next_state = 2000;  end 
1444: begin if(four_bit_hash == 0) next_state = 1445; else  next_state = 2000;  end 
1445: begin if(four_bit_hash == 0) next_state = 1446; else  next_state = 2000;  end 
1446: begin if(four_bit_hash == 0) next_state = 1447; else  next_state = 2000;  end 
1447: begin if(four_bit_hash == 0) next_state = 1448; else  next_state = 2000;  end 
1448: begin if(four_bit_hash == 0) next_state = 1449; else  next_state = 2000;  end 
1449: begin if(four_bit_hash == 0) next_state = 1450; else  next_state = 2000;  end 
1450: begin if(four_bit_hash == 0) next_state = 1451; else  next_state = 2000;  end 
1451: begin if(four_bit_hash == 0) next_state = 1452; else  next_state = 2000;  end 
1452: begin if(four_bit_hash == 0) next_state = 1453; else  next_state = 2000;  end 
1453: begin if(four_bit_hash == 0) next_state = 1454; else  next_state = 2000;  end 
1454: begin if(four_bit_hash == 0) next_state = 1455; else  next_state = 2000;  end 
1455: begin if(four_bit_hash == 0) next_state = 1456; else  next_state = 2000;  end 
1456: begin if(four_bit_hash == 0) next_state = 1457; else  next_state = 2000;  end 
1457: begin if(four_bit_hash == 0) next_state = 1458; else  next_state = 2000;  end 
1458: begin if(four_bit_hash == 0) next_state = 1459; else  next_state = 2000;  end 
1459: begin if(four_bit_hash == 0) next_state = 1460; else  next_state = 2000;  end 
1460: begin if(four_bit_hash == 0) next_state = 1461; else  next_state = 2000;  end 
1461: begin if(four_bit_hash == 0) next_state = 1462; else  next_state = 2000;  end 
1462: begin if(four_bit_hash == 0) next_state = 1463; else  next_state = 2000;  end 
1463: begin if(four_bit_hash == 0) next_state = 1464; else  next_state = 2000;  end 
1464: begin if(four_bit_hash == 0) next_state = 1465; else  next_state = 2000;  end 
1465: begin if(four_bit_hash == 0) next_state = 1466; else  next_state = 2000;  end 
1466: begin if(four_bit_hash == 0) next_state = 1467; else  next_state = 2000;  end 
1467: begin if(four_bit_hash == 0) next_state = 1468; else  next_state = 2000;  end 
1468: begin if(four_bit_hash == 0) next_state = 1469; else  next_state = 2000;  end 
1469: begin if(four_bit_hash == 0) next_state = 1470; else  next_state = 2000;  end 
1470: begin if(four_bit_hash == 0) next_state = 1471; else  next_state = 2000;  end 
1471: begin if(four_bit_hash == 0) next_state = 1472; else  next_state = 2000;  end 
1472: begin if(four_bit_hash == 0) next_state = 1473; else  next_state = 2000;  end 
1473: begin if(four_bit_hash == 0) next_state = 1474; else  next_state = 2000;  end 
1474: begin if(four_bit_hash == 0) next_state = 1475; else  next_state = 2000;  end 
1475: begin if(four_bit_hash == 0) next_state = 1476; else  next_state = 2000;  end 
1476: begin if(four_bit_hash == 0) next_state = 1477; else  next_state = 2000;  end 
1477: begin if(four_bit_hash == 0) next_state = 1478; else  next_state = 2000;  end 
1478: begin if(four_bit_hash == 0) next_state = 1479; else  next_state = 2000;  end 
1479: begin if(four_bit_hash == 0) next_state = 1480; else  next_state = 2000;  end 
1480: begin if(four_bit_hash == 0) next_state = 1481; else  next_state = 2000;  end 
1481: begin if(four_bit_hash == 0) next_state = 1482; else  next_state = 2000;  end 
1482: begin if(four_bit_hash == 0) next_state = 1483; else  next_state = 2000;  end 
1483: begin if(four_bit_hash == 0) next_state = 1484; else  next_state = 2000;  end 
1484: begin if(four_bit_hash == 0) next_state = 1485; else  next_state = 2000;  end 
1485: begin if(four_bit_hash == 0) next_state = 1486; else  next_state = 2000;  end 
1486: begin if(four_bit_hash == 0) next_state = 1487; else  next_state = 2000;  end 
1487: begin if(four_bit_hash == 0) next_state = 1488; else  next_state = 2000;  end 
1488: begin if(four_bit_hash == 0) next_state = 1489; else  next_state = 2000;  end 
1489: begin if(four_bit_hash == 0) next_state = 1490; else  next_state = 2000;  end 
1490: begin if(four_bit_hash == 0) next_state = 1491; else  next_state = 2000;  end 
1491: begin if(four_bit_hash == 0) next_state = 1492; else  next_state = 2000;  end 
1492: begin if(four_bit_hash == 0) next_state = 1493; else  next_state = 2000;  end 
1493: begin if(four_bit_hash == 0) next_state = 1494; else  next_state = 2000;  end 
1494: begin if(four_bit_hash == 0) next_state = 1495; else  next_state = 2000;  end 
1495: begin if(four_bit_hash == 0) next_state = 1496; else  next_state = 2000;  end 
1496: begin if(four_bit_hash == 0) next_state = 1497; else  next_state = 2000;  end 
1497: begin if(four_bit_hash == 0) next_state = 1498; else  next_state = 2000;  end 
1498: begin if(four_bit_hash == 0) next_state = 1499; else  next_state = 2000;  end 
1499: begin if(four_bit_hash == 0) next_state = 1500; else  next_state = 2000;  end 
1500: begin if(four_bit_hash == 0) next_state = 1501; else  next_state = 2000;  end 
1501: begin if(four_bit_hash == 0) next_state = 1502; else  next_state = 2000;  end 
1502: begin if(four_bit_hash == 0) next_state = 1503; else  next_state = 2000;  end 
1503: begin if(four_bit_hash == 0) next_state = 1504; else  next_state = 2000;  end 
1504: begin if(four_bit_hash == 0) next_state = 1505; else  next_state = 2000;  end 
1505: begin if(four_bit_hash == 0) next_state = 1506; else  next_state = 2000;  end 
1506: begin if(four_bit_hash == 0) next_state = 1507; else  next_state = 2000;  end 
1507: begin if(four_bit_hash == 0) next_state = 1508; else  next_state = 2000;  end 
1508: begin if(four_bit_hash == 0) next_state = 1509; else  next_state = 2000;  end 
1509: begin if(four_bit_hash == 0) next_state = 1510; else  next_state = 2000;  end 
1510: begin if(four_bit_hash == 0) next_state = 1511; else  next_state = 2000;  end 
1511: begin if(four_bit_hash == 0) next_state = 1512; else  next_state = 2000;  end 
1512: begin if(four_bit_hash == 0) next_state = 1513; else  next_state = 2000;  end 
1513: begin if(four_bit_hash == 0) next_state = 1514; else  next_state = 2000;  end 
1514: begin if(four_bit_hash == 0) next_state = 1515; else  next_state = 2000;  end 
1515: begin if(four_bit_hash == 0) next_state = 1516; else  next_state = 2000;  end 
1516: begin if(four_bit_hash == 0) next_state = 1517; else  next_state = 2000;  end 
1517: begin if(four_bit_hash == 0) next_state = 1518; else  next_state = 2000;  end 
1518: begin if(four_bit_hash == 0) next_state = 1519; else  next_state = 2000;  end 
1519: begin if(four_bit_hash == 0) next_state = 1520; else  next_state = 2000;  end 
1520: begin if(four_bit_hash == 0) next_state = 1521; else  next_state = 2000;  end 
1521: begin if(four_bit_hash == 0) next_state = 1522; else  next_state = 2000;  end 
1522: begin if(four_bit_hash == 0) next_state = 1523; else  next_state = 2000;  end 
1523: begin if(four_bit_hash == 0) next_state = 1524; else  next_state = 2000;  end 
1524: begin if(four_bit_hash == 0) next_state = 1525; else  next_state = 2000;  end 
1525: begin if(four_bit_hash == 0) next_state = 1526; else  next_state = 2000;  end 
1526: begin if(four_bit_hash == 0) next_state = 1527; else  next_state = 2000;  end 
1527: begin if(four_bit_hash == 0) next_state = 1528; else  next_state = 2000;  end 
1528: begin if(four_bit_hash == 0) next_state = 1529; else  next_state = 2000;  end 
1529: begin if(four_bit_hash == 0) next_state = 1530; else  next_state = 2000;  end 
1530: begin if(four_bit_hash == 0) next_state = 1531; else  next_state = 2000;  end 
1531: begin if(four_bit_hash == 0) next_state = 1532; else  next_state = 2000;  end 
1532: begin if(four_bit_hash == 0) next_state = 1533; else  next_state = 2000;  end 
1533: begin if(four_bit_hash == 0) next_state = 1534; else  next_state = 2000;  end 
1534: begin if(four_bit_hash == 0) next_state = 1535; else  next_state = 2000;  end 
1535: begin if(four_bit_hash == 0) next_state = 1536; else  next_state = 2000;  end 
1536: begin if(four_bit_hash == 0) next_state = 1537; else  next_state = 2000;  end 
1537: begin if(four_bit_hash == 0) next_state = 1538; else  next_state = 2000;  end 
1538: begin if(four_bit_hash == 0) next_state = 1539; else  next_state = 2000;  end 
1539: begin if(four_bit_hash == 0) next_state = 1540; else  next_state = 2000;  end 
1540: begin if(four_bit_hash == 0) next_state = 1541; else  next_state = 2000;  end 
1541: begin if(four_bit_hash == 0) next_state = 1542; else  next_state = 2000;  end 
1542: begin if(four_bit_hash == 0) next_state = 1543; else  next_state = 2000;  end 
1543: begin if(four_bit_hash == 0) next_state = 1544; else  next_state = 2000;  end 
1544: begin if(four_bit_hash == 0) next_state = 1545; else  next_state = 2000;  end 
1545: begin if(four_bit_hash == 0) next_state = 1546; else  next_state = 2000;  end 
1546: begin if(four_bit_hash == 0) next_state = 1547; else  next_state = 2000;  end 
1547: begin if(four_bit_hash == 0) next_state = 1548; else  next_state = 2000;  end 
1548: begin if(four_bit_hash == 0) next_state = 1549; else  next_state = 2000;  end 
1549: begin if(four_bit_hash == 0) next_state = 1550; else  next_state = 2000;  end 
1550: begin if(four_bit_hash == 0) next_state = 1551; else  next_state = 2000;  end 
1551: begin if(four_bit_hash == 0) next_state = 1552; else  next_state = 2000;  end 
1552: begin if(four_bit_hash == 0) next_state = 1553; else  next_state = 2000;  end  
2000: begin packet_drop_signal_register  = 1'b1; end
default: begin next_state = 0;end
endcase
end

assign packet_drop_signal =packet_drop_signal_out;
endmodule