library verilog;
use verilog.vl_types.all;
entity user_data_path is
    generic(
        DATA_WIDTH      : integer := 64;
        CTRL_WIDTH      : vl_notype;
        UDP_REG_SRC_WIDTH: integer := 2;
        NUM_OUTPUT_QUEUES: integer := 8;
        NUM_INPUT_QUEUES: integer := 8;
        SRAM_DATA_WIDTH : vl_notype;
        SRAM_ADDR_WIDTH : integer := 19
    );
    port(
        in_data_0       : in     vl_logic_vector;
        in_ctrl_0       : in     vl_logic_vector;
        in_wr_0         : in     vl_logic;
        in_rdy_0        : out    vl_logic;
        in_data_1       : in     vl_logic_vector;
        in_ctrl_1       : in     vl_logic_vector;
        in_wr_1         : in     vl_logic;
        in_rdy_1        : out    vl_logic;
        in_data_2       : in     vl_logic_vector;
        in_ctrl_2       : in     vl_logic_vector;
        in_wr_2         : in     vl_logic;
        in_rdy_2        : out    vl_logic;
        in_data_3       : in     vl_logic_vector;
        in_ctrl_3       : in     vl_logic_vector;
        in_wr_3         : in     vl_logic;
        in_rdy_3        : out    vl_logic;
        in_data_4       : in     vl_logic_vector;
        in_ctrl_4       : in     vl_logic_vector;
        in_wr_4         : in     vl_logic;
        in_rdy_4        : out    vl_logic;
        in_data_5       : in     vl_logic_vector;
        in_ctrl_5       : in     vl_logic_vector;
        in_wr_5         : in     vl_logic;
        in_rdy_5        : out    vl_logic;
        in_data_6       : in     vl_logic_vector;
        in_ctrl_6       : in     vl_logic_vector;
        in_wr_6         : in     vl_logic;
        in_rdy_6        : out    vl_logic;
        in_data_7       : in     vl_logic_vector;
        in_ctrl_7       : in     vl_logic_vector;
        in_wr_7         : in     vl_logic;
        in_rdy_7        : out    vl_logic;
        out_data_0      : out    vl_logic_vector;
        out_ctrl_0      : out    vl_logic_vector;
        out_wr_0        : out    vl_logic;
        out_rdy_0       : in     vl_logic;
        out_data_1      : out    vl_logic_vector;
        out_ctrl_1      : out    vl_logic_vector;
        out_wr_1        : out    vl_logic;
        out_rdy_1       : in     vl_logic;
        out_data_2      : out    vl_logic_vector;
        out_ctrl_2      : out    vl_logic_vector;
        out_wr_2        : out    vl_logic;
        out_rdy_2       : in     vl_logic;
        out_data_3      : out    vl_logic_vector;
        out_ctrl_3      : out    vl_logic_vector;
        out_wr_3        : out    vl_logic;
        out_rdy_3       : in     vl_logic;
        out_data_4      : out    vl_logic_vector;
        out_ctrl_4      : out    vl_logic_vector;
        out_wr_4        : out    vl_logic;
        out_rdy_4       : in     vl_logic;
        out_data_5      : out    vl_logic_vector;
        out_ctrl_5      : out    vl_logic_vector;
        out_wr_5        : out    vl_logic;
        out_rdy_5       : in     vl_logic;
        out_data_6      : out    vl_logic_vector;
        out_ctrl_6      : out    vl_logic_vector;
        out_wr_6        : out    vl_logic;
        out_rdy_6       : in     vl_logic;
        out_data_7      : out    vl_logic_vector;
        out_ctrl_7      : out    vl_logic_vector;
        out_wr_7        : out    vl_logic;
        out_rdy_7       : in     vl_logic;
        wr_0_addr       : out    vl_logic_vector;
        wr_0_req        : out    vl_logic;
        wr_0_ack        : in     vl_logic;
        wr_0_data       : out    vl_logic_vector;
        rd_0_ack        : in     vl_logic;
        rd_0_data       : in     vl_logic_vector;
        rd_0_vld        : in     vl_logic;
        rd_0_addr       : out    vl_logic_vector;
        rd_0_req        : out    vl_logic;
        reg_req         : in     vl_logic;
        reg_ack         : out    vl_logic;
        reg_rd_wr_L     : in     vl_logic;
        reg_addr        : in     vl_logic_vector(22 downto 0);
        reg_rd_data     : out    vl_logic_vector(31 downto 0);
        reg_wr_data     : in     vl_logic_vector(31 downto 0);
        reset           : in     vl_logic;
        clk             : in     vl_logic;
        statemac_clk    : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CTRL_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of UDP_REG_SRC_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_OUTPUT_QUEUES : constant is 1;
    attribute mti_svvh_generic_type of NUM_INPUT_QUEUES : constant is 1;
    attribute mti_svvh_generic_type of SRAM_DATA_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of SRAM_ADDR_WIDTH : constant is 1;
end user_data_path;
