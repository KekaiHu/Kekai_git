library verilog;
use verilog.vl_types.all;
entity oq_regs_ctrl is
    generic(
        SRAM_ADDR_WIDTH : integer := 13;
        CTRL_WIDTH      : integer := 8;
        NUM_OUTPUT_QUEUES: integer := 8;
        NUM_OQ_WIDTH    : vl_notype;
        NUM_REGS_USED   : integer := 17;
        ADDR_WIDTH      : vl_notype;
        MAX_PKT         : vl_notype;
        MIN_PKT         : vl_notype;
        PKTS_IN_RAM_WIDTH: vl_notype;
        PKT_LEN_WIDTH   : integer := 11;
        PKT_WORDS_WIDTH : vl_notype
    );
    port(
        enable          : out    vl_logic_vector;
        reg_req         : in     vl_logic;
        reg_rd_wr_L_held: in     vl_logic;
        reg_data_held   : in     vl_logic_vector(31 downto 0);
        addr            : in     vl_logic_vector;
        q_addr          : in     vl_logic_vector;
        result_ready    : out    vl_logic;
        reg_result      : out    vl_logic_vector(31 downto 0);
        initialize      : out    vl_logic;
        initialize_oq   : out    vl_logic_vector;
        reg_addr        : out    vl_logic_vector;
        num_pkt_bytes_stored_reg_req: out    vl_logic;
        num_pkt_bytes_stored_reg_ack: in     vl_logic;
        num_pkt_bytes_stored_reg_wr: out    vl_logic;
        num_pkt_bytes_stored_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkt_bytes_stored_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_overhead_bytes_stored_reg_req: out    vl_logic;
        num_overhead_bytes_stored_reg_ack: in     vl_logic;
        num_overhead_bytes_stored_reg_wr: out    vl_logic;
        num_overhead_bytes_stored_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_overhead_bytes_stored_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_pkts_stored_reg_req: out    vl_logic;
        num_pkts_stored_reg_ack: in     vl_logic;
        num_pkts_stored_reg_wr: out    vl_logic;
        num_pkts_stored_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkts_stored_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_pkts_dropped_reg_req: out    vl_logic;
        num_pkts_dropped_reg_ack: in     vl_logic;
        num_pkts_dropped_reg_wr: out    vl_logic;
        num_pkts_dropped_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkts_dropped_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_pkt_bytes_removed_reg_req: out    vl_logic;
        num_pkt_bytes_removed_reg_ack: in     vl_logic;
        num_pkt_bytes_removed_reg_wr: out    vl_logic;
        num_pkt_bytes_removed_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkt_bytes_removed_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_overhead_bytes_removed_reg_req: out    vl_logic;
        num_overhead_bytes_removed_reg_ack: in     vl_logic;
        num_overhead_bytes_removed_reg_wr: out    vl_logic;
        num_overhead_bytes_removed_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_overhead_bytes_removed_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_pkts_removed_reg_req: out    vl_logic;
        num_pkts_removed_reg_ack: in     vl_logic;
        num_pkts_removed_reg_wr: out    vl_logic;
        num_pkts_removed_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkts_removed_reg_rd_data: in     vl_logic_vector(31 downto 0);
        oq_addr_hi_reg_req: out    vl_logic;
        oq_addr_hi_reg_ack: in     vl_logic;
        oq_addr_hi_reg_wr: out    vl_logic;
        oq_addr_hi_reg_wr_data: out    vl_logic_vector(31 downto 0);
        oq_addr_hi_reg_rd_data: in     vl_logic_vector(31 downto 0);
        oq_addr_lo_reg_req: out    vl_logic;
        oq_addr_lo_reg_ack: in     vl_logic;
        oq_addr_lo_reg_wr: out    vl_logic;
        oq_addr_lo_reg_wr_data: out    vl_logic_vector(31 downto 0);
        oq_addr_lo_reg_rd_data: in     vl_logic_vector(31 downto 0);
        oq_wr_addr_reg_req: out    vl_logic;
        oq_wr_addr_reg_ack: in     vl_logic;
        oq_wr_addr_reg_wr: out    vl_logic;
        oq_wr_addr_reg_wr_data: out    vl_logic_vector(31 downto 0);
        oq_wr_addr_reg_rd_data: in     vl_logic_vector(31 downto 0);
        oq_rd_addr_reg_req: out    vl_logic;
        oq_rd_addr_reg_ack: in     vl_logic;
        oq_rd_addr_reg_wr: out    vl_logic;
        oq_rd_addr_reg_wr_data: out    vl_logic_vector(31 downto 0);
        oq_rd_addr_reg_rd_data: in     vl_logic_vector(31 downto 0);
        max_pkts_in_q_reg_req: out    vl_logic;
        max_pkts_in_q_reg_ack: in     vl_logic;
        max_pkts_in_q_reg_wr: out    vl_logic;
        max_pkts_in_q_reg_wr_data: out    vl_logic_vector(31 downto 0);
        max_pkts_in_q_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_pkts_in_q_reg_req: out    vl_logic;
        num_pkts_in_q_reg_ack: in     vl_logic;
        num_pkts_in_q_reg_wr: out    vl_logic;
        num_pkts_in_q_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_pkts_in_q_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_words_left_reg_req: out    vl_logic;
        num_words_left_reg_ack: in     vl_logic;
        num_words_left_reg_wr: out    vl_logic;
        num_words_left_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_words_left_reg_rd_data: in     vl_logic_vector(31 downto 0);
        num_words_in_q_reg_req: out    vl_logic;
        num_words_in_q_reg_ack: in     vl_logic;
        num_words_in_q_reg_wr: out    vl_logic;
        num_words_in_q_reg_wr_data: out    vl_logic_vector(31 downto 0);
        num_words_in_q_reg_rd_data: in     vl_logic_vector(31 downto 0);
        oq_full_thresh_reg_req: out    vl_logic;
        oq_full_thresh_reg_ack: in     vl_logic;
        oq_full_thresh_reg_wr: out    vl_logic;
        oq_full_thresh_reg_wr_data: out    vl_logic_vector(31 downto 0);
        oq_full_thresh_reg_rd_data: in     vl_logic_vector(31 downto 0);
        clk             : in     vl_logic;
        reset           : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SRAM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of CTRL_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of NUM_OUTPUT_QUEUES : constant is 1;
    attribute mti_svvh_generic_type of NUM_OQ_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of NUM_REGS_USED : constant is 1;
    attribute mti_svvh_generic_type of ADDR_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of MAX_PKT : constant is 3;
    attribute mti_svvh_generic_type of MIN_PKT : constant is 3;
    attribute mti_svvh_generic_type of PKTS_IN_RAM_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of PKT_LEN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of PKT_WORDS_WIDTH : constant is 3;
end oq_regs_ctrl;
